------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80d0f80c",
3 => x"3a0b0b80",
4 => x"c8d40400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d0",
162 => x"94738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d0f40c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c7e23f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"90822d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8ed02d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80e0e4",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80e0",
307 => x"e4085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480d0",
314 => x"f408802e",
315 => x"a43880d0",
316 => x"f808822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80e0e40c",
320 => x"82a0800b",
321 => x"80e0e80c",
322 => x"8290800b",
323 => x"80e0ec0c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80e0e4",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"e0e80cf8",
330 => x"80808480",
331 => x"0b80e0ec",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80e0",
335 => x"e40c80c0",
336 => x"a880940b",
337 => x"80e0e80c",
338 => x"80d0a40b",
339 => x"80e0ec0c",
340 => x"04ff3d0d",
341 => x"80e0f033",
342 => x"5170a738",
343 => x"80d18008",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"d1800c70",
348 => x"2d80d180",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80e0",
352 => x"f034833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80e0e008",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"e0e0510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404803d",
366 => x"0d80e0fc",
367 => x"08811180",
368 => x"e0fc0c51",
369 => x"823d0d04",
370 => x"f73d0d7b",
371 => x"54870b89",
372 => x"3d80d184",
373 => x"08585855",
374 => x"7417748f",
375 => x"06175353",
376 => x"71337334",
377 => x"73842aff",
378 => x"16565474",
379 => x"8025e938",
380 => x"800b8b3d",
381 => x"34765188",
382 => x"ae3f8b3d",
383 => x"0d04e93d",
384 => x"0d80e0fc",
385 => x"08973d95",
386 => x"3d933d91",
387 => x"3d80e0fc",
388 => x"08575c5c",
389 => x"5c5c5c7b",
390 => x"722e828f",
391 => x"3880d0bc",
392 => x"5188843f",
393 => x"80e0fc08",
394 => x"8c808008",
395 => x"8c808408",
396 => x"80d0cc54",
397 => x"59545c87",
398 => x"ee3f7254",
399 => x"870b80d1",
400 => x"84085755",
401 => x"741b748f",
402 => x"06175353",
403 => x"71337334",
404 => x"73842aff",
405 => x"16565474",
406 => x"8025e938",
407 => x"800b993d",
408 => x"347a5187",
409 => x"c23f80d0",
410 => x"d05187bb",
411 => x"3f765487",
412 => x"0b80d184",
413 => x"08575574",
414 => x"1a748f06",
415 => x"17545772",
416 => x"33773473",
417 => x"842aff16",
418 => x"56547480",
419 => x"25e93880",
420 => x"0b963d34",
421 => x"7951878f",
422 => x"3ff8bb95",
423 => x"86a10b8c",
424 => x"80800c81",
425 => x"91d1acf8",
426 => x"0b8c8084",
427 => x"0c8c8080",
428 => x"088c8084",
429 => x"0880d0cc",
430 => x"53585586",
431 => x"ea3f7454",
432 => x"870b80d1",
433 => x"84085755",
434 => x"7419748f",
435 => x"06175353",
436 => x"71337334",
437 => x"73842aff",
438 => x"16565474",
439 => x"8025e938",
440 => x"800b933d",
441 => x"34785186",
442 => x"be3f80d0",
443 => x"d05186b7",
444 => x"3f765487",
445 => x"0b80d184",
446 => x"08575574",
447 => x"18748f06",
448 => x"17545772",
449 => x"33773473",
450 => x"842aff16",
451 => x"56547480",
452 => x"25e93880",
453 => x"0b903d34",
454 => x"7751868b",
455 => x"3f80e0fc",
456 => x"08527b72",
457 => x"2e098106",
458 => x"fdf33880",
459 => x"d0d45185",
460 => x"f63f8c80",
461 => x"80088c80",
462 => x"840880d0",
463 => x"cc535853",
464 => x"85e53f72",
465 => x"54870b80",
466 => x"d1840857",
467 => x"55fdf539",
468 => x"bc0802bc",
469 => x"0cf93d0d",
470 => x"800bbc08",
471 => x"fc050cbc",
472 => x"08880508",
473 => x"8025ab38",
474 => x"bc088805",
475 => x"0830bc08",
476 => x"88050c80",
477 => x"0bbc08f4",
478 => x"050cbc08",
479 => x"fc050888",
480 => x"38810bbc",
481 => x"08f4050c",
482 => x"bc08f405",
483 => x"08bc08fc",
484 => x"050cbc08",
485 => x"8c050880",
486 => x"25ab38bc",
487 => x"088c0508",
488 => x"30bc088c",
489 => x"050c800b",
490 => x"bc08f005",
491 => x"0cbc08fc",
492 => x"05088838",
493 => x"810bbc08",
494 => x"f0050cbc",
495 => x"08f00508",
496 => x"bc08fc05",
497 => x"0c8053bc",
498 => x"088c0508",
499 => x"52bc0888",
500 => x"05085181",
501 => x"a73fb008",
502 => x"70bc08f8",
503 => x"050c54bc",
504 => x"08fc0508",
505 => x"802e8c38",
506 => x"bc08f805",
507 => x"0830bc08",
508 => x"f8050cbc",
509 => x"08f80508",
510 => x"70b00c54",
511 => x"893d0dbc",
512 => x"0c04bc08",
513 => x"02bc0cfb",
514 => x"3d0d800b",
515 => x"bc08fc05",
516 => x"0cbc0888",
517 => x"05088025",
518 => x"9338bc08",
519 => x"88050830",
520 => x"bc088805",
521 => x"0c810bbc",
522 => x"08fc050c",
523 => x"bc088c05",
524 => x"0880258c",
525 => x"38bc088c",
526 => x"050830bc",
527 => x"088c050c",
528 => x"8153bc08",
529 => x"8c050852",
530 => x"bc088805",
531 => x"0851ad3f",
532 => x"b00870bc",
533 => x"08f8050c",
534 => x"54bc08fc",
535 => x"0508802e",
536 => x"8c38bc08",
537 => x"f8050830",
538 => x"bc08f805",
539 => x"0cbc08f8",
540 => x"050870b0",
541 => x"0c54873d",
542 => x"0dbc0c04",
543 => x"bc0802bc",
544 => x"0cfd3d0d",
545 => x"810bbc08",
546 => x"fc050c80",
547 => x"0bbc08f8",
548 => x"050cbc08",
549 => x"8c0508bc",
550 => x"08880508",
551 => x"27ac38bc",
552 => x"08fc0508",
553 => x"802ea338",
554 => x"800bbc08",
555 => x"8c050824",
556 => x"9938bc08",
557 => x"8c050810",
558 => x"bc088c05",
559 => x"0cbc08fc",
560 => x"050810bc",
561 => x"08fc050c",
562 => x"c939bc08",
563 => x"fc050880",
564 => x"2e80c938",
565 => x"bc088c05",
566 => x"08bc0888",
567 => x"050826a1",
568 => x"38bc0888",
569 => x"0508bc08",
570 => x"8c050831",
571 => x"bc088805",
572 => x"0cbc08f8",
573 => x"0508bc08",
574 => x"fc050807",
575 => x"bc08f805",
576 => x"0cbc08fc",
577 => x"0508812a",
578 => x"bc08fc05",
579 => x"0cbc088c",
580 => x"0508812a",
581 => x"bc088c05",
582 => x"0cffaf39",
583 => x"bc089005",
584 => x"08802e8f",
585 => x"38bc0888",
586 => x"050870bc",
587 => x"08f4050c",
588 => x"518d39bc",
589 => x"08f80508",
590 => x"70bc08f4",
591 => x"050c51bc",
592 => x"08f40508",
593 => x"b00c853d",
594 => x"0dbc0c04",
595 => x"fc3d0d76",
596 => x"70797b55",
597 => x"5555558f",
598 => x"72278c38",
599 => x"72750783",
600 => x"06517080",
601 => x"2ea738ff",
602 => x"125271ff",
603 => x"2e983872",
604 => x"70810554",
605 => x"33747081",
606 => x"055634ff",
607 => x"125271ff",
608 => x"2e098106",
609 => x"ea3874b0",
610 => x"0c863d0d",
611 => x"04745172",
612 => x"70840554",
613 => x"08717084",
614 => x"05530c72",
615 => x"70840554",
616 => x"08717084",
617 => x"05530c72",
618 => x"70840554",
619 => x"08717084",
620 => x"05530c72",
621 => x"70840554",
622 => x"08717084",
623 => x"05530cf0",
624 => x"1252718f",
625 => x"26c93883",
626 => x"72279538",
627 => x"72708405",
628 => x"54087170",
629 => x"8405530c",
630 => x"fc125271",
631 => x"8326ed38",
632 => x"7054ff83",
633 => x"39f73d0d",
634 => x"7c705253",
635 => x"80ca3f72",
636 => x"54b00855",
637 => x"0b0b80d0",
638 => x"e0568157",
639 => x"b0088105",
640 => x"5a8b3de4",
641 => x"11595382",
642 => x"59f41352",
643 => x"7b881108",
644 => x"52538183",
645 => x"3fb00830",
646 => x"70b00807",
647 => x"9f2c8a07",
648 => x"b00c538b",
649 => x"3d0d04ff",
650 => x"3d0d7352",
651 => x"80d18808",
652 => x"51ffb23f",
653 => x"833d0d04",
654 => x"fd3d0d75",
655 => x"70718306",
656 => x"53555270",
657 => x"b8387170",
658 => x"087009f7",
659 => x"fbfdff12",
660 => x"0670f884",
661 => x"82818006",
662 => x"51515253",
663 => x"709d3884",
664 => x"13700870",
665 => x"09f7fbfd",
666 => x"ff120670",
667 => x"f8848281",
668 => x"80065151",
669 => x"52537080",
670 => x"2ee53872",
671 => x"52713351",
672 => x"70802e8a",
673 => x"38811270",
674 => x"33525270",
675 => x"f8387174",
676 => x"31b00c85",
677 => x"3d0d04f2",
678 => x"3d0d6062",
679 => x"88110870",
680 => x"57575f5a",
681 => x"74802e81",
682 => x"8f388c1a",
683 => x"2270832a",
684 => x"81327081",
685 => x"06515558",
686 => x"73863890",
687 => x"1a089138",
688 => x"795190a1",
689 => x"3fff54b0",
690 => x"0880ed38",
691 => x"8c1a2258",
692 => x"7d085780",
693 => x"7883ffff",
694 => x"0670812a",
695 => x"70810651",
696 => x"56575573",
697 => x"752e80d7",
698 => x"38749038",
699 => x"76088418",
700 => x"08881959",
701 => x"56597480",
702 => x"2ef23874",
703 => x"54888075",
704 => x"27843888",
705 => x"80547353",
706 => x"78529c1a",
707 => x"0851a41a",
708 => x"0854732d",
709 => x"800bb008",
710 => x"2582e638",
711 => x"b0081975",
712 => x"b008317f",
713 => x"880508b0",
714 => x"08317061",
715 => x"88050c56",
716 => x"565973ff",
717 => x"b4388054",
718 => x"73b00c90",
719 => x"3d0d0475",
720 => x"81327081",
721 => x"06764151",
722 => x"5473802e",
723 => x"81c13874",
724 => x"90387608",
725 => x"84180888",
726 => x"19595659",
727 => x"74802ef2",
728 => x"38881a08",
729 => x"7883ffff",
730 => x"0670892a",
731 => x"70810651",
732 => x"56595673",
733 => x"802e82fa",
734 => x"38757527",
735 => x"8d387787",
736 => x"2a708106",
737 => x"51547382",
738 => x"b5387476",
739 => x"27833874",
740 => x"56755378",
741 => x"52790851",
742 => x"85823f88",
743 => x"1a087631",
744 => x"881b0c79",
745 => x"08167a0c",
746 => x"74567519",
747 => x"7577317f",
748 => x"88050878",
749 => x"31706188",
750 => x"050c5656",
751 => x"5973802e",
752 => x"fef4388c",
753 => x"1a2258ff",
754 => x"86397778",
755 => x"5479537b",
756 => x"525684c8",
757 => x"3f881a08",
758 => x"7831881b",
759 => x"0c790818",
760 => x"7a0c7c76",
761 => x"315d7c8e",
762 => x"3879518f",
763 => x"db3fb008",
764 => x"818f38b0",
765 => x"085f7519",
766 => x"7577317f",
767 => x"88050878",
768 => x"31706188",
769 => x"050c5656",
770 => x"5973802e",
771 => x"fea83874",
772 => x"81833876",
773 => x"08841808",
774 => x"88195956",
775 => x"5974802e",
776 => x"f2387453",
777 => x"8a527851",
778 => x"82d33fb0",
779 => x"08793181",
780 => x"055db008",
781 => x"84388115",
782 => x"5d815f7c",
783 => x"58747d27",
784 => x"83387458",
785 => x"941a0888",
786 => x"1b081157",
787 => x"5c807a08",
788 => x"5c54901a",
789 => x"087b2783",
790 => x"38815475",
791 => x"78258438",
792 => x"73ba387b",
793 => x"7824fee2",
794 => x"387b5378",
795 => x"529c1a08",
796 => x"51a41a08",
797 => x"54732db0",
798 => x"0856b008",
799 => x"8024fee2",
800 => x"388c1a22",
801 => x"80c00754",
802 => x"738c1b23",
803 => x"ff5473b0",
804 => x"0c903d0d",
805 => x"047effa3",
806 => x"38ff8739",
807 => x"75537852",
808 => x"7a5182f8",
809 => x"3f790816",
810 => x"7a0c7951",
811 => x"8e9a3fb0",
812 => x"08cf387c",
813 => x"76315d7c",
814 => x"febc38fe",
815 => x"ac39901a",
816 => x"087a0871",
817 => x"31761170",
818 => x"565a5752",
819 => x"80d18808",
820 => x"51848c3f",
821 => x"b008802e",
822 => x"ffa738b0",
823 => x"08901b0c",
824 => x"b008167a",
825 => x"0c77941b",
826 => x"0c74881b",
827 => x"0c7456fd",
828 => x"99397908",
829 => x"58901a08",
830 => x"78278338",
831 => x"81547575",
832 => x"27843873",
833 => x"b338941a",
834 => x"08567575",
835 => x"2680d338",
836 => x"75537852",
837 => x"9c1a0851",
838 => x"a41a0854",
839 => x"732db008",
840 => x"56b00880",
841 => x"24fd8338",
842 => x"8c1a2280",
843 => x"c0075473",
844 => x"8c1b23ff",
845 => x"54fed739",
846 => x"75537852",
847 => x"775181dc",
848 => x"3f790816",
849 => x"7a0c7951",
850 => x"8cfe3fb0",
851 => x"08802efc",
852 => x"d9388c1a",
853 => x"2280c007",
854 => x"54738c1b",
855 => x"23ff54fe",
856 => x"ad397475",
857 => x"54795378",
858 => x"525681b0",
859 => x"3f881a08",
860 => x"7531881b",
861 => x"0c790815",
862 => x"7a0cfcae",
863 => x"39fa3d0d",
864 => x"7a790288",
865 => x"05a70533",
866 => x"56525383",
867 => x"73278a38",
868 => x"70830652",
869 => x"71802ea8",
870 => x"38ff1353",
871 => x"72ff2e97",
872 => x"38703352",
873 => x"73722e91",
874 => x"388111ff",
875 => x"14545172",
876 => x"ff2e0981",
877 => x"06eb3880",
878 => x"5170b00c",
879 => x"883d0d04",
880 => x"70725755",
881 => x"83517582",
882 => x"802914ff",
883 => x"12525670",
884 => x"8025f338",
885 => x"837327bf",
886 => x"38740876",
887 => x"327009f7",
888 => x"fbfdff12",
889 => x"0670f884",
890 => x"82818006",
891 => x"51515170",
892 => x"802e9938",
893 => x"74518052",
894 => x"70335773",
895 => x"772effb9",
896 => x"38811181",
897 => x"13535183",
898 => x"7227ed38",
899 => x"fc138416",
900 => x"56537283",
901 => x"26c33874",
902 => x"51fefe39",
903 => x"fa3d0d78",
904 => x"7a7c7272",
905 => x"72575757",
906 => x"59565674",
907 => x"7627b238",
908 => x"76155175",
909 => x"7127aa38",
910 => x"707717ff",
911 => x"14545553",
912 => x"71ff2e96",
913 => x"38ff14ff",
914 => x"14545472",
915 => x"337434ff",
916 => x"125271ff",
917 => x"2e098106",
918 => x"ec3875b0",
919 => x"0c883d0d",
920 => x"04768f26",
921 => x"9738ff12",
922 => x"5271ff2e",
923 => x"ed387270",
924 => x"81055433",
925 => x"74708105",
926 => x"5634eb39",
927 => x"74760783",
928 => x"065170e2",
929 => x"38757554",
930 => x"51727084",
931 => x"05540871",
932 => x"70840553",
933 => x"0c727084",
934 => x"05540871",
935 => x"70840553",
936 => x"0c727084",
937 => x"05540871",
938 => x"70840553",
939 => x"0c727084",
940 => x"05540871",
941 => x"70840553",
942 => x"0cf01252",
943 => x"718f26c9",
944 => x"38837227",
945 => x"95387270",
946 => x"84055408",
947 => x"71708405",
948 => x"530cfc12",
949 => x"52718326",
950 => x"ed387054",
951 => x"ff8839ef",
952 => x"3d0d6365",
953 => x"67405d42",
954 => x"7b802e84",
955 => x"fa386151",
956 => x"a5b43ff8",
957 => x"1c708412",
958 => x"0870fc06",
959 => x"70628b05",
960 => x"70f80641",
961 => x"59455b5c",
962 => x"41579674",
963 => x"2782c338",
964 => x"807b247e",
965 => x"7c260759",
966 => x"80547874",
967 => x"2e098106",
968 => x"82a93877",
969 => x"7b2581fc",
970 => x"38771780",
971 => x"d8c40b88",
972 => x"05085e56",
973 => x"7c762e84",
974 => x"bd388416",
975 => x"0870fe06",
976 => x"17841108",
977 => x"81065155",
978 => x"5573828b",
979 => x"3874fc06",
980 => x"597c762e",
981 => x"84dd3877",
982 => x"195f7e7b",
983 => x"2581fd38",
984 => x"79810654",
985 => x"7382bf38",
986 => x"76770831",
987 => x"841108fc",
988 => x"06565a75",
989 => x"802e9138",
990 => x"7c762e84",
991 => x"ea387419",
992 => x"1859787b",
993 => x"25848938",
994 => x"79802e82",
995 => x"99387715",
996 => x"567a7624",
997 => x"8290388c",
998 => x"1a08881b",
999 => x"08718c12",
1000 => x"0c88120c",
1001 => x"55797659",
1002 => x"57881761",
1003 => x"fc055759",
1004 => x"75a42685",
1005 => x"ef387b79",
1006 => x"55559376",
1007 => x"2780c938",
1008 => x"7b708405",
1009 => x"5d087c56",
1010 => x"790c7470",
1011 => x"84055608",
1012 => x"8c180c90",
1013 => x"17549b76",
1014 => x"27ae3874",
1015 => x"70840556",
1016 => x"08740c74",
1017 => x"70840556",
1018 => x"0894180c",
1019 => x"981754a3",
1020 => x"76279538",
1021 => x"74708405",
1022 => x"5608740c",
1023 => x"74708405",
1024 => x"56089c18",
1025 => x"0ca01754",
1026 => x"74708405",
1027 => x"56087470",
1028 => x"8405560c",
1029 => x"74708405",
1030 => x"56087470",
1031 => x"8405560c",
1032 => x"7408740c",
1033 => x"777b3156",
1034 => x"758f2680",
1035 => x"c9388417",
1036 => x"08810678",
1037 => x"0784180c",
1038 => x"77178411",
1039 => x"08810784",
1040 => x"120c5461",
1041 => x"51a2e03f",
1042 => x"88175473",
1043 => x"b00c933d",
1044 => x"0d04905b",
1045 => x"fdba3978",
1046 => x"56fe8539",
1047 => x"8c160888",
1048 => x"1708718c",
1049 => x"120c8812",
1050 => x"0c557e70",
1051 => x"7c315758",
1052 => x"8f7627ff",
1053 => x"b9387a17",
1054 => x"84180881",
1055 => x"067c0784",
1056 => x"190c7681",
1057 => x"0784120c",
1058 => x"76118411",
1059 => x"08810784",
1060 => x"120c5588",
1061 => x"05526151",
1062 => x"8cf63f61",
1063 => x"51a2883f",
1064 => x"881754ff",
1065 => x"a6397d52",
1066 => x"615194f5",
1067 => x"3fb00859",
1068 => x"b008802e",
1069 => x"81a338b0",
1070 => x"08f80560",
1071 => x"840508fe",
1072 => x"06610555",
1073 => x"5776742e",
1074 => x"83e638fc",
1075 => x"185675a4",
1076 => x"2681aa38",
1077 => x"7bb00855",
1078 => x"55937627",
1079 => x"80d83874",
1080 => x"70840556",
1081 => x"08b00870",
1082 => x"8405b00c",
1083 => x"0cb00875",
1084 => x"70840557",
1085 => x"08717084",
1086 => x"05530c54",
1087 => x"9b7627b6",
1088 => x"38747084",
1089 => x"05560874",
1090 => x"70840556",
1091 => x"0c747084",
1092 => x"05560874",
1093 => x"70840556",
1094 => x"0ca37627",
1095 => x"99387470",
1096 => x"84055608",
1097 => x"74708405",
1098 => x"560c7470",
1099 => x"84055608",
1100 => x"74708405",
1101 => x"560c7470",
1102 => x"84055608",
1103 => x"74708405",
1104 => x"560c7470",
1105 => x"84055608",
1106 => x"74708405",
1107 => x"560c7408",
1108 => x"740c7b52",
1109 => x"61518bb8",
1110 => x"3f6151a0",
1111 => x"ca3f7854",
1112 => x"73b00c93",
1113 => x"3d0d047d",
1114 => x"52615193",
1115 => x"b43fb008",
1116 => x"b00c933d",
1117 => x"0d048416",
1118 => x"0855fbd1",
1119 => x"3975537b",
1120 => x"52b00851",
1121 => x"efc63f7b",
1122 => x"5261518b",
1123 => x"833fca39",
1124 => x"8c160888",
1125 => x"1708718c",
1126 => x"120c8812",
1127 => x"0c558c1a",
1128 => x"08881b08",
1129 => x"718c120c",
1130 => x"88120c55",
1131 => x"79795957",
1132 => x"fbf73977",
1133 => x"19901c55",
1134 => x"55737524",
1135 => x"fba2387a",
1136 => x"177080d8",
1137 => x"c40b8805",
1138 => x"0c757c31",
1139 => x"81078412",
1140 => x"0c5d8417",
1141 => x"0881067b",
1142 => x"0784180c",
1143 => x"61519fc7",
1144 => x"3f881754",
1145 => x"fce53974",
1146 => x"1918901c",
1147 => x"555d737d",
1148 => x"24fb9538",
1149 => x"8c1a0888",
1150 => x"1b08718c",
1151 => x"120c8812",
1152 => x"0c55881a",
1153 => x"61fc0557",
1154 => x"5975a426",
1155 => x"81ae387b",
1156 => x"79555593",
1157 => x"762780c9",
1158 => x"387b7084",
1159 => x"055d087c",
1160 => x"56790c74",
1161 => x"70840556",
1162 => x"088c1b0c",
1163 => x"901a549b",
1164 => x"7627ae38",
1165 => x"74708405",
1166 => x"5608740c",
1167 => x"74708405",
1168 => x"5608941b",
1169 => x"0c981a54",
1170 => x"a3762795",
1171 => x"38747084",
1172 => x"05560874",
1173 => x"0c747084",
1174 => x"0556089c",
1175 => x"1b0ca01a",
1176 => x"54747084",
1177 => x"05560874",
1178 => x"70840556",
1179 => x"0c747084",
1180 => x"05560874",
1181 => x"70840556",
1182 => x"0c740874",
1183 => x"0c7a1a70",
1184 => x"80d8c40b",
1185 => x"88050c7d",
1186 => x"7c318107",
1187 => x"84120c54",
1188 => x"841a0881",
1189 => x"067b0784",
1190 => x"1b0c6151",
1191 => x"9e893f78",
1192 => x"54fdbd39",
1193 => x"75537b52",
1194 => x"7851eda0",
1195 => x"3ffaf539",
1196 => x"841708fc",
1197 => x"06186058",
1198 => x"58fae939",
1199 => x"75537b52",
1200 => x"7851ed88",
1201 => x"3f7a1a70",
1202 => x"80d8c40b",
1203 => x"88050c7d",
1204 => x"7c318107",
1205 => x"84120c54",
1206 => x"841a0881",
1207 => x"067b0784",
1208 => x"1b0cffb6",
1209 => x"39fa3d0d",
1210 => x"7880d188",
1211 => x"085455b8",
1212 => x"1308802e",
1213 => x"81b5388c",
1214 => x"15227083",
1215 => x"ffff0670",
1216 => x"832a8132",
1217 => x"70810651",
1218 => x"55555672",
1219 => x"802e80dc",
1220 => x"3873842a",
1221 => x"81328106",
1222 => x"57ff5376",
1223 => x"80f63873",
1224 => x"822a7081",
1225 => x"06515372",
1226 => x"802eb938",
1227 => x"b0150854",
1228 => x"73802e9c",
1229 => x"3880c015",
1230 => x"5373732e",
1231 => x"8f387352",
1232 => x"80d18808",
1233 => x"5187c93f",
1234 => x"8c152256",
1235 => x"76b0160c",
1236 => x"75db0653",
1237 => x"728c1623",
1238 => x"800b8416",
1239 => x"0c901508",
1240 => x"750c7256",
1241 => x"75880753",
1242 => x"728c1623",
1243 => x"90150880",
1244 => x"2e80c038",
1245 => x"8c152270",
1246 => x"81065553",
1247 => x"739d3872",
1248 => x"812a7081",
1249 => x"06515372",
1250 => x"85389415",
1251 => x"08547388",
1252 => x"160c8053",
1253 => x"72b00c88",
1254 => x"3d0d0480",
1255 => x"0b88160c",
1256 => x"94150830",
1257 => x"98160c80",
1258 => x"53ea3972",
1259 => x"5182fb3f",
1260 => x"fec53974",
1261 => x"518ce83f",
1262 => x"8c152270",
1263 => x"81065553",
1264 => x"73802eff",
1265 => x"ba38d439",
1266 => x"f83d0d7a",
1267 => x"5877802e",
1268 => x"81993880",
1269 => x"d1880854",
1270 => x"b8140880",
1271 => x"2e80ed38",
1272 => x"8c182270",
1273 => x"902b7090",
1274 => x"2c70832a",
1275 => x"81328106",
1276 => x"5c515754",
1277 => x"7880cd38",
1278 => x"90180857",
1279 => x"76802e80",
1280 => x"c3387708",
1281 => x"77317779",
1282 => x"0c768306",
1283 => x"7a585555",
1284 => x"73853894",
1285 => x"18085675",
1286 => x"88190c80",
1287 => x"7525a538",
1288 => x"74537652",
1289 => x"9c180851",
1290 => x"a4180854",
1291 => x"732d800b",
1292 => x"b0082580",
1293 => x"c938b008",
1294 => x"1775b008",
1295 => x"31565774",
1296 => x"8024dd38",
1297 => x"800bb00c",
1298 => x"8a3d0d04",
1299 => x"735181da",
1300 => x"3f8c1822",
1301 => x"70902b70",
1302 => x"902c7083",
1303 => x"2a813281",
1304 => x"065c5157",
1305 => x"5478dd38",
1306 => x"ff8e39a7",
1307 => x"c85280d1",
1308 => x"88085189",
1309 => x"f13fb008",
1310 => x"b00c8a3d",
1311 => x"0d048c18",
1312 => x"2280c007",
1313 => x"54738c19",
1314 => x"23ff0bb0",
1315 => x"0c8a3d0d",
1316 => x"04803d0d",
1317 => x"72518071",
1318 => x"0c800b84",
1319 => x"120c800b",
1320 => x"88120c02",
1321 => x"8e05228c",
1322 => x"12230292",
1323 => x"05228e12",
1324 => x"23800b90",
1325 => x"120c800b",
1326 => x"94120c80",
1327 => x"0b98120c",
1328 => x"709c120c",
1329 => x"80c3dc0b",
1330 => x"a0120c80",
1331 => x"c4a80ba4",
1332 => x"120c80c5",
1333 => x"a40ba812",
1334 => x"0c80c5f5",
1335 => x"0bac120c",
1336 => x"823d0d04",
1337 => x"fa3d0d79",
1338 => x"7080dc29",
1339 => x"8c11547a",
1340 => x"5356578c",
1341 => x"ac3fb008",
1342 => x"b0085556",
1343 => x"b008802e",
1344 => x"a238b008",
1345 => x"8c055480",
1346 => x"0bb0080c",
1347 => x"76b00884",
1348 => x"050c73b0",
1349 => x"0888050c",
1350 => x"74538052",
1351 => x"735197f7",
1352 => x"3f755473",
1353 => x"b00c883d",
1354 => x"0d04fc3d",
1355 => x"0d76acbd",
1356 => x"0bbc120c",
1357 => x"55810bb8",
1358 => x"160c800b",
1359 => x"84dc160c",
1360 => x"830b84e0",
1361 => x"160c84e8",
1362 => x"1584e416",
1363 => x"0c745480",
1364 => x"53845284",
1365 => x"150851fe",
1366 => x"b83f7454",
1367 => x"81538952",
1368 => x"88150851",
1369 => x"feab3f74",
1370 => x"5482538a",
1371 => x"528c1508",
1372 => x"51fe9e3f",
1373 => x"863d0d04",
1374 => x"f93d0d79",
1375 => x"80d18808",
1376 => x"5457b813",
1377 => x"08802e80",
1378 => x"c83884dc",
1379 => x"13568816",
1380 => x"08841708",
1381 => x"ff055555",
1382 => x"8074249f",
1383 => x"388c1522",
1384 => x"70902b70",
1385 => x"902c5154",
1386 => x"5872802e",
1387 => x"80ca3880",
1388 => x"dc15ff15",
1389 => x"55557380",
1390 => x"25e33875",
1391 => x"08537280",
1392 => x"2e9f3872",
1393 => x"56881608",
1394 => x"841708ff",
1395 => x"055555c8",
1396 => x"397251fe",
1397 => x"d53f80d1",
1398 => x"880884dc",
1399 => x"0556ffae",
1400 => x"39845276",
1401 => x"51fdfd3f",
1402 => x"b008760c",
1403 => x"b008802e",
1404 => x"80c038b0",
1405 => x"0856ce39",
1406 => x"810b8c16",
1407 => x"2372750c",
1408 => x"7288160c",
1409 => x"7284160c",
1410 => x"7290160c",
1411 => x"7294160c",
1412 => x"7298160c",
1413 => x"ff0b8e16",
1414 => x"2372b016",
1415 => x"0c72b416",
1416 => x"0c7280c4",
1417 => x"160c7280",
1418 => x"c8160c74",
1419 => x"b00c893d",
1420 => x"0d048c77",
1421 => x"0c800bb0",
1422 => x"0c893d0d",
1423 => x"04ff3d0d",
1424 => x"a7c85273",
1425 => x"51869f3f",
1426 => x"833d0d04",
1427 => x"803d0d80",
1428 => x"d1880851",
1429 => x"e83f823d",
1430 => x"0d04fb3d",
1431 => x"0d777052",
1432 => x"5696c33f",
1433 => x"80d8c40b",
1434 => x"88050884",
1435 => x"1108fc06",
1436 => x"707b319f",
1437 => x"ef05e080",
1438 => x"06e08005",
1439 => x"565653a0",
1440 => x"80742494",
1441 => x"38805275",
1442 => x"51969d3f",
1443 => x"80d8cc08",
1444 => x"155372b0",
1445 => x"082e8f38",
1446 => x"7551968b",
1447 => x"3f805372",
1448 => x"b00c873d",
1449 => x"0d047330",
1450 => x"52755195",
1451 => x"fb3fb008",
1452 => x"ff2ea838",
1453 => x"80d8c40b",
1454 => x"88050875",
1455 => x"75318107",
1456 => x"84120c53",
1457 => x"80d88808",
1458 => x"743180d8",
1459 => x"880c7551",
1460 => x"95d53f81",
1461 => x"0bb00c87",
1462 => x"3d0d0480",
1463 => x"52755195",
1464 => x"c73f80d8",
1465 => x"c40b8805",
1466 => x"08b00871",
1467 => x"3156538f",
1468 => x"7525ffa4",
1469 => x"38b00880",
1470 => x"d8b80831",
1471 => x"80d8880c",
1472 => x"74810784",
1473 => x"140c7551",
1474 => x"959d3f80",
1475 => x"53ff9039",
1476 => x"f63d0d7c",
1477 => x"7e545b72",
1478 => x"802e8283",
1479 => x"387a5195",
1480 => x"853ff813",
1481 => x"84110870",
1482 => x"fe067013",
1483 => x"841108fc",
1484 => x"065d5859",
1485 => x"545880d8",
1486 => x"cc08752e",
1487 => x"82de3878",
1488 => x"84160c80",
1489 => x"73810654",
1490 => x"5a727a2e",
1491 => x"81d53878",
1492 => x"15841108",
1493 => x"81065153",
1494 => x"72a03878",
1495 => x"17577981",
1496 => x"e6388815",
1497 => x"08537280",
1498 => x"d8cc2e82",
1499 => x"f9388c15",
1500 => x"08708c15",
1501 => x"0c738812",
1502 => x"0c567681",
1503 => x"0784190c",
1504 => x"76187771",
1505 => x"0c537981",
1506 => x"913883ff",
1507 => x"772781c8",
1508 => x"3876892a",
1509 => x"77832a56",
1510 => x"5372802e",
1511 => x"bf387686",
1512 => x"2ab80555",
1513 => x"847327b4",
1514 => x"3880db13",
1515 => x"55947327",
1516 => x"ab38768c",
1517 => x"2a80ee05",
1518 => x"5580d473",
1519 => x"279e3876",
1520 => x"8f2a80f7",
1521 => x"055582d4",
1522 => x"73279138",
1523 => x"76922a80",
1524 => x"fc05558a",
1525 => x"d4732784",
1526 => x"3880fe55",
1527 => x"74101010",
1528 => x"80d8c405",
1529 => x"88110855",
1530 => x"5673762e",
1531 => x"82b33884",
1532 => x"1408fc06",
1533 => x"53767327",
1534 => x"8d388814",
1535 => x"08547376",
1536 => x"2e098106",
1537 => x"ea388c14",
1538 => x"08708c1a",
1539 => x"0c74881a",
1540 => x"0c788812",
1541 => x"0c56778c",
1542 => x"150c7a51",
1543 => x"93893f8c",
1544 => x"3d0d0477",
1545 => x"08787131",
1546 => x"59770588",
1547 => x"19085457",
1548 => x"7280d8cc",
1549 => x"2e80e038",
1550 => x"8c180870",
1551 => x"8c150c73",
1552 => x"88120c56",
1553 => x"fe893988",
1554 => x"15088c16",
1555 => x"08708c13",
1556 => x"0c578817",
1557 => x"0cfea339",
1558 => x"76832a70",
1559 => x"54558075",
1560 => x"24819838",
1561 => x"72822c81",
1562 => x"712b80d8",
1563 => x"c8080780",
1564 => x"d8c40b84",
1565 => x"050c5374",
1566 => x"10101080",
1567 => x"d8c40588",
1568 => x"11085556",
1569 => x"758c190c",
1570 => x"7388190c",
1571 => x"7788170c",
1572 => x"778c150c",
1573 => x"ff843981",
1574 => x"5afdb439",
1575 => x"78177381",
1576 => x"06545772",
1577 => x"98387708",
1578 => x"78713159",
1579 => x"77058c19",
1580 => x"08881a08",
1581 => x"718c120c",
1582 => x"88120c57",
1583 => x"57768107",
1584 => x"84190c77",
1585 => x"80d8c40b",
1586 => x"88050c80",
1587 => x"d8c00877",
1588 => x"26fec738",
1589 => x"80d8bc08",
1590 => x"527a51fa",
1591 => x"fd3f7a51",
1592 => x"91c53ffe",
1593 => x"ba398178",
1594 => x"8c150c78",
1595 => x"88150c73",
1596 => x"8c1a0c73",
1597 => x"881a0c5a",
1598 => x"fd803983",
1599 => x"1570822c",
1600 => x"81712b80",
1601 => x"d8c80807",
1602 => x"80d8c40b",
1603 => x"84050c51",
1604 => x"53741010",
1605 => x"1080d8c4",
1606 => x"05881108",
1607 => x"5556fee4",
1608 => x"39745380",
1609 => x"7524a738",
1610 => x"72822c81",
1611 => x"712b80d8",
1612 => x"c8080780",
1613 => x"d8c40b84",
1614 => x"050c5375",
1615 => x"8c190c73",
1616 => x"88190c77",
1617 => x"88170c77",
1618 => x"8c150cfd",
1619 => x"cd398315",
1620 => x"70822c81",
1621 => x"712b80d8",
1622 => x"c8080780",
1623 => x"d8c40b84",
1624 => x"050c5153",
1625 => x"d639f93d",
1626 => x"0d797b58",
1627 => x"53800b80",
1628 => x"d1880853",
1629 => x"5672722e",
1630 => x"80c03884",
1631 => x"dc135574",
1632 => x"762eb738",
1633 => x"88150884",
1634 => x"1608ff05",
1635 => x"54548073",
1636 => x"249d388c",
1637 => x"14227090",
1638 => x"2b70902c",
1639 => x"51535871",
1640 => x"80d83880",
1641 => x"dc14ff14",
1642 => x"54547280",
1643 => x"25e53874",
1644 => x"085574d0",
1645 => x"3880d188",
1646 => x"085284dc",
1647 => x"12557480",
1648 => x"2eb13888",
1649 => x"15088416",
1650 => x"08ff0554",
1651 => x"54807324",
1652 => x"9c388c14",
1653 => x"2270902b",
1654 => x"70902c51",
1655 => x"535871ad",
1656 => x"3880dc14",
1657 => x"ff145454",
1658 => x"728025e6",
1659 => x"38740855",
1660 => x"74d13875",
1661 => x"b00c893d",
1662 => x"0d047351",
1663 => x"762d75b0",
1664 => x"080780dc",
1665 => x"15ff1555",
1666 => x"5556ff9e",
1667 => x"39735176",
1668 => x"2d75b008",
1669 => x"0780dc15",
1670 => x"ff155555",
1671 => x"56ca39ea",
1672 => x"3d0d688c",
1673 => x"11227081",
1674 => x"2a810657",
1675 => x"58567480",
1676 => x"e4388e16",
1677 => x"2270902b",
1678 => x"70902c51",
1679 => x"55588074",
1680 => x"24b13898",
1681 => x"3dc40553",
1682 => x"735280d1",
1683 => x"88085192",
1684 => x"ac3f800b",
1685 => x"b0082497",
1686 => x"387983e0",
1687 => x"80065473",
1688 => x"80c0802e",
1689 => x"818f3873",
1690 => x"8280802e",
1691 => x"8191388c",
1692 => x"16225776",
1693 => x"90800754",
1694 => x"738c1723",
1695 => x"88805280",
1696 => x"d1880851",
1697 => x"819b3fb0",
1698 => x"089d388c",
1699 => x"16228207",
1700 => x"54738c17",
1701 => x"2380c316",
1702 => x"70770c90",
1703 => x"170c810b",
1704 => x"94170c98",
1705 => x"3d0d0480",
1706 => x"d18808ac",
1707 => x"bd0bbc12",
1708 => x"0c548c16",
1709 => x"22818007",
1710 => x"54738c17",
1711 => x"23b00876",
1712 => x"0cb00890",
1713 => x"170c8880",
1714 => x"0b94170c",
1715 => x"74802ed3",
1716 => x"388e1622",
1717 => x"70902b70",
1718 => x"902c5355",
1719 => x"5898ae3f",
1720 => x"b008802e",
1721 => x"ffbd388c",
1722 => x"16228107",
1723 => x"54738c17",
1724 => x"23983d0d",
1725 => x"04810b8c",
1726 => x"17225855",
1727 => x"fef539a8",
1728 => x"160880c5",
1729 => x"a42e0981",
1730 => x"06fee438",
1731 => x"8c162288",
1732 => x"80075473",
1733 => x"8c172388",
1734 => x"800b80cc",
1735 => x"170cfedc",
1736 => x"39f33d0d",
1737 => x"7f618b11",
1738 => x"70f8065c",
1739 => x"55555e72",
1740 => x"96268338",
1741 => x"90598079",
1742 => x"24747a26",
1743 => x"07538054",
1744 => x"72742e09",
1745 => x"810680cb",
1746 => x"387d518c",
1747 => x"d93f7883",
1748 => x"f72680c6",
1749 => x"3878832a",
1750 => x"70101010",
1751 => x"80d8c405",
1752 => x"8c110859",
1753 => x"595a7678",
1754 => x"2e83b038",
1755 => x"841708fc",
1756 => x"06568c17",
1757 => x"08881808",
1758 => x"718c120c",
1759 => x"88120c58",
1760 => x"75178411",
1761 => x"08810784",
1762 => x"120c537d",
1763 => x"518c983f",
1764 => x"88175473",
1765 => x"b00c8f3d",
1766 => x"0d047889",
1767 => x"2a79832a",
1768 => x"5b537280",
1769 => x"2ebf3878",
1770 => x"862ab805",
1771 => x"5a847327",
1772 => x"b43880db",
1773 => x"135a9473",
1774 => x"27ab3878",
1775 => x"8c2a80ee",
1776 => x"055a80d4",
1777 => x"73279e38",
1778 => x"788f2a80",
1779 => x"f7055a82",
1780 => x"d4732791",
1781 => x"3878922a",
1782 => x"80fc055a",
1783 => x"8ad47327",
1784 => x"843880fe",
1785 => x"5a791010",
1786 => x"1080d8c4",
1787 => x"058c1108",
1788 => x"58557675",
1789 => x"2ea33884",
1790 => x"1708fc06",
1791 => x"707a3155",
1792 => x"56738f24",
1793 => x"88d53873",
1794 => x"8025fee6",
1795 => x"388c1708",
1796 => x"5776752e",
1797 => x"098106df",
1798 => x"38811a5a",
1799 => x"80d8d408",
1800 => x"577680d8",
1801 => x"cc2e82c0",
1802 => x"38841708",
1803 => x"fc06707a",
1804 => x"31555673",
1805 => x"8f2481f9",
1806 => x"3880d8cc",
1807 => x"0b80d8d8",
1808 => x"0c80d8cc",
1809 => x"0b80d8d4",
1810 => x"0c738025",
1811 => x"feb23883",
1812 => x"ff762783",
1813 => x"df387589",
1814 => x"2a76832a",
1815 => x"55537280",
1816 => x"2ebf3875",
1817 => x"862ab805",
1818 => x"54847327",
1819 => x"b43880db",
1820 => x"13549473",
1821 => x"27ab3875",
1822 => x"8c2a80ee",
1823 => x"055480d4",
1824 => x"73279e38",
1825 => x"758f2a80",
1826 => x"f7055482",
1827 => x"d4732791",
1828 => x"3875922a",
1829 => x"80fc0554",
1830 => x"8ad47327",
1831 => x"843880fe",
1832 => x"54731010",
1833 => x"1080d8c4",
1834 => x"05881108",
1835 => x"56587478",
1836 => x"2e86cf38",
1837 => x"841508fc",
1838 => x"06537573",
1839 => x"278d3888",
1840 => x"15085574",
1841 => x"782e0981",
1842 => x"06ea388c",
1843 => x"150880d8",
1844 => x"c40b8405",
1845 => x"08718c1a",
1846 => x"0c76881a",
1847 => x"0c788813",
1848 => x"0c788c18",
1849 => x"0c5d5879",
1850 => x"53807a24",
1851 => x"83e63872",
1852 => x"822c8171",
1853 => x"2b5c537a",
1854 => x"7c268198",
1855 => x"387b7b06",
1856 => x"537282f1",
1857 => x"3879fc06",
1858 => x"84055a7a",
1859 => x"10707d06",
1860 => x"545b7282",
1861 => x"e038841a",
1862 => x"5af13988",
1863 => x"178c1108",
1864 => x"58587678",
1865 => x"2e098106",
1866 => x"fcc23882",
1867 => x"1a5afdec",
1868 => x"39781779",
1869 => x"81078419",
1870 => x"0c7080d8",
1871 => x"d80c7080",
1872 => x"d8d40c80",
1873 => x"d8cc0b8c",
1874 => x"120c8c11",
1875 => x"0888120c",
1876 => x"74810784",
1877 => x"120c7411",
1878 => x"75710c51",
1879 => x"537d5188",
1880 => x"c63f8817",
1881 => x"54fcac39",
1882 => x"80d8c40b",
1883 => x"8405087a",
1884 => x"545c7980",
1885 => x"25fef838",
1886 => x"82da397a",
1887 => x"097c0670",
1888 => x"80d8c40b",
1889 => x"84050c5c",
1890 => x"7a105b7a",
1891 => x"7c268538",
1892 => x"7a85b838",
1893 => x"80d8c40b",
1894 => x"88050870",
1895 => x"841208fc",
1896 => x"06707c31",
1897 => x"7c72268f",
1898 => x"72250757",
1899 => x"575c5d55",
1900 => x"72802e80",
1901 => x"db38797a",
1902 => x"1680d8bc",
1903 => x"081b9011",
1904 => x"5a55575b",
1905 => x"80d8b808",
1906 => x"ff2e8838",
1907 => x"a08f13e0",
1908 => x"80065776",
1909 => x"527d5187",
1910 => x"cf3fb008",
1911 => x"54b008ff",
1912 => x"2e9038b0",
1913 => x"08762782",
1914 => x"99387480",
1915 => x"d8c42e82",
1916 => x"913880d8",
1917 => x"c40b8805",
1918 => x"08558415",
1919 => x"08fc0670",
1920 => x"7a317a72",
1921 => x"268f7225",
1922 => x"07525553",
1923 => x"7283e638",
1924 => x"74798107",
1925 => x"84170c79",
1926 => x"167080d8",
1927 => x"c40b8805",
1928 => x"0c758107",
1929 => x"84120c54",
1930 => x"7e525786",
1931 => x"fa3f8817",
1932 => x"54fae039",
1933 => x"75832a70",
1934 => x"54548074",
1935 => x"24819b38",
1936 => x"72822c81",
1937 => x"712b80d8",
1938 => x"c8080770",
1939 => x"80d8c40b",
1940 => x"84050c75",
1941 => x"10101080",
1942 => x"d8c40588",
1943 => x"1108585a",
1944 => x"5d53778c",
1945 => x"180c7488",
1946 => x"180c7688",
1947 => x"190c768c",
1948 => x"160cfcf3",
1949 => x"39797a10",
1950 => x"101080d8",
1951 => x"c4057057",
1952 => x"595d8c15",
1953 => x"08577675",
1954 => x"2ea33884",
1955 => x"1708fc06",
1956 => x"707a3155",
1957 => x"56738f24",
1958 => x"83ca3873",
1959 => x"80258481",
1960 => x"388c1708",
1961 => x"5776752e",
1962 => x"098106df",
1963 => x"38881581",
1964 => x"1b708306",
1965 => x"555b5572",
1966 => x"c9387c83",
1967 => x"06537280",
1968 => x"2efdb838",
1969 => x"ff1df819",
1970 => x"595d8818",
1971 => x"08782eea",
1972 => x"38fdb539",
1973 => x"831a53fc",
1974 => x"96398314",
1975 => x"70822c81",
1976 => x"712b80d8",
1977 => x"c8080770",
1978 => x"80d8c40b",
1979 => x"84050c76",
1980 => x"10101080",
1981 => x"d8c40588",
1982 => x"1108595b",
1983 => x"5e5153fe",
1984 => x"e13980d8",
1985 => x"88081758",
1986 => x"b008762e",
1987 => x"818d3880",
1988 => x"d8b808ff",
1989 => x"2e83ec38",
1990 => x"73763118",
1991 => x"80d8880c",
1992 => x"73870670",
1993 => x"57537280",
1994 => x"2e883888",
1995 => x"73317015",
1996 => x"55567614",
1997 => x"9fff06a0",
1998 => x"80713117",
1999 => x"70547f53",
2000 => x"575384e4",
2001 => x"3fb00853",
2002 => x"b008ff2e",
2003 => x"81a03880",
2004 => x"d8880816",
2005 => x"7080d888",
2006 => x"0c747580",
2007 => x"d8c40b88",
2008 => x"050c7476",
2009 => x"31187081",
2010 => x"07515556",
2011 => x"587b80d8",
2012 => x"c42e839c",
2013 => x"38798f26",
2014 => x"82cb3881",
2015 => x"0b84150c",
2016 => x"841508fc",
2017 => x"06707a31",
2018 => x"7a72268f",
2019 => x"72250752",
2020 => x"55537280",
2021 => x"2efcf938",
2022 => x"80db39b0",
2023 => x"089fff06",
2024 => x"5372feeb",
2025 => x"387780d8",
2026 => x"880c80d8",
2027 => x"c40b8805",
2028 => x"087b1881",
2029 => x"0784120c",
2030 => x"5580d8b4",
2031 => x"08782786",
2032 => x"387780d8",
2033 => x"b40c80d8",
2034 => x"b0087827",
2035 => x"fcac3877",
2036 => x"80d8b00c",
2037 => x"841508fc",
2038 => x"06707a31",
2039 => x"7a72268f",
2040 => x"72250752",
2041 => x"55537280",
2042 => x"2efca538",
2043 => x"88398074",
2044 => x"5456fedb",
2045 => x"397d5183",
2046 => x"ae3f800b",
2047 => x"b00c8f3d",
2048 => x"0d047353",
2049 => x"807424a9",
2050 => x"3872822c",
2051 => x"81712b80",
2052 => x"d8c80807",
2053 => x"7080d8c4",
2054 => x"0b84050c",
2055 => x"5d53778c",
2056 => x"180c7488",
2057 => x"180c7688",
2058 => x"190c768c",
2059 => x"160cf9b7",
2060 => x"39831470",
2061 => x"822c8171",
2062 => x"2b80d8c8",
2063 => x"08077080",
2064 => x"d8c40b84",
2065 => x"050c5e51",
2066 => x"53d4397b",
2067 => x"7b065372",
2068 => x"fca33884",
2069 => x"1a7b105c",
2070 => x"5af139ff",
2071 => x"1a811151",
2072 => x"5af7b939",
2073 => x"78177981",
2074 => x"0784190c",
2075 => x"8c180888",
2076 => x"1908718c",
2077 => x"120c8812",
2078 => x"0c597080",
2079 => x"d8d80c70",
2080 => x"80d8d40c",
2081 => x"80d8cc0b",
2082 => x"8c120c8c",
2083 => x"11088812",
2084 => x"0c748107",
2085 => x"84120c74",
2086 => x"1175710c",
2087 => x"5153f9bd",
2088 => x"39751784",
2089 => x"11088107",
2090 => x"84120c53",
2091 => x"8c170888",
2092 => x"1808718c",
2093 => x"120c8812",
2094 => x"0c587d51",
2095 => x"81e93f88",
2096 => x"1754f5cf",
2097 => x"39728415",
2098 => x"0cf41af8",
2099 => x"0670841e",
2100 => x"08810607",
2101 => x"841e0c70",
2102 => x"1d545b85",
2103 => x"0b84140c",
2104 => x"850b8814",
2105 => x"0c8f7b27",
2106 => x"fdcf3888",
2107 => x"1c527d51",
2108 => x"ec9e3f80",
2109 => x"d8c40b88",
2110 => x"050880d8",
2111 => x"88085955",
2112 => x"fdb73977",
2113 => x"80d8880c",
2114 => x"7380d8b8",
2115 => x"0cfc9139",
2116 => x"7284150c",
2117 => x"fda339fc",
2118 => x"3d0d7679",
2119 => x"71028c05",
2120 => x"9f053357",
2121 => x"55535583",
2122 => x"72278a38",
2123 => x"74830651",
2124 => x"70802ea2",
2125 => x"38ff1252",
2126 => x"71ff2e93",
2127 => x"38737370",
2128 => x"81055534",
2129 => x"ff125271",
2130 => x"ff2e0981",
2131 => x"06ef3874",
2132 => x"b00c863d",
2133 => x"0d047474",
2134 => x"882b7507",
2135 => x"7071902b",
2136 => x"07515451",
2137 => x"8f7227a5",
2138 => x"38727170",
2139 => x"8405530c",
2140 => x"72717084",
2141 => x"05530c72",
2142 => x"71708405",
2143 => x"530c7271",
2144 => x"70840553",
2145 => x"0cf01252",
2146 => x"718f26dd",
2147 => x"38837227",
2148 => x"90387271",
2149 => x"70840553",
2150 => x"0cfc1252",
2151 => x"718326f2",
2152 => x"387053ff",
2153 => x"90390404",
2154 => x"fd3d0d80",
2155 => x"0b80e180",
2156 => x"0c765184",
2157 => x"ee3fb008",
2158 => x"53b008ff",
2159 => x"2e883872",
2160 => x"b00c853d",
2161 => x"0d0480e1",
2162 => x"80085473",
2163 => x"802ef038",
2164 => x"7574710c",
2165 => x"5272b00c",
2166 => x"853d0d04",
2167 => x"f93d0d79",
2168 => x"7c557b54",
2169 => x"8e112270",
2170 => x"902b7090",
2171 => x"2c555780",
2172 => x"d1880853",
2173 => x"585683f3",
2174 => x"3fb00857",
2175 => x"800bb008",
2176 => x"24933880",
2177 => x"d01608b0",
2178 => x"080580d0",
2179 => x"170c76b0",
2180 => x"0c893d0d",
2181 => x"048c1622",
2182 => x"83dfff06",
2183 => x"55748c17",
2184 => x"2376b00c",
2185 => x"893d0d04",
2186 => x"fa3d0d78",
2187 => x"8c112270",
2188 => x"882a7081",
2189 => x"06515758",
2190 => x"5674a938",
2191 => x"8c162283",
2192 => x"dfff0655",
2193 => x"748c1723",
2194 => x"7a547953",
2195 => x"8e162270",
2196 => x"902b7090",
2197 => x"2c545680",
2198 => x"d1880852",
2199 => x"5681b23f",
2200 => x"883d0d04",
2201 => x"82548053",
2202 => x"8e162270",
2203 => x"902b7090",
2204 => x"2c545680",
2205 => x"d1880852",
2206 => x"5782b83f",
2207 => x"8c162283",
2208 => x"dfff0655",
2209 => x"748c1723",
2210 => x"7a547953",
2211 => x"8e162270",
2212 => x"902b7090",
2213 => x"2c545680",
2214 => x"d1880852",
2215 => x"5680f23f",
2216 => x"883d0d04",
2217 => x"f93d0d79",
2218 => x"7c557b54",
2219 => x"8e112270",
2220 => x"902b7090",
2221 => x"2c555780",
2222 => x"d1880853",
2223 => x"585681f3",
2224 => x"3fb00857",
2225 => x"b008ff2e",
2226 => x"99388c16",
2227 => x"22a08007",
2228 => x"55748c17",
2229 => x"23b00880",
2230 => x"d0170c76",
2231 => x"b00c893d",
2232 => x"0d048c16",
2233 => x"2283dfff",
2234 => x"0655748c",
2235 => x"172376b0",
2236 => x"0c893d0d",
2237 => x"04fe3d0d",
2238 => x"748e1122",
2239 => x"70902b70",
2240 => x"902c5551",
2241 => x"515380d1",
2242 => x"880851bd",
2243 => x"3f843d0d",
2244 => x"04fb3d0d",
2245 => x"800b80e1",
2246 => x"800c7a53",
2247 => x"79527851",
2248 => x"82fb3fb0",
2249 => x"0855b008",
2250 => x"ff2e8838",
2251 => x"74b00c87",
2252 => x"3d0d0480",
2253 => x"e1800856",
2254 => x"75802ef0",
2255 => x"38777671",
2256 => x"0c5474b0",
2257 => x"0c873d0d",
2258 => x"04fd3d0d",
2259 => x"800b80e1",
2260 => x"800c7651",
2261 => x"84d03fb0",
2262 => x"0853b008",
2263 => x"ff2e8838",
2264 => x"72b00c85",
2265 => x"3d0d0480",
2266 => x"e1800854",
2267 => x"73802ef0",
2268 => x"38757471",
2269 => x"0c5272b0",
2270 => x"0c853d0d",
2271 => x"04fc3d0d",
2272 => x"800b80e1",
2273 => x"800c7852",
2274 => x"775186b8",
2275 => x"3fb00854",
2276 => x"b008ff2e",
2277 => x"883873b0",
2278 => x"0c863d0d",
2279 => x"0480e180",
2280 => x"08557480",
2281 => x"2ef03876",
2282 => x"75710c53",
2283 => x"73b00c86",
2284 => x"3d0d04fb",
2285 => x"3d0d800b",
2286 => x"80e1800c",
2287 => x"7a537952",
2288 => x"78518494",
2289 => x"3fb00855",
2290 => x"b008ff2e",
2291 => x"883874b0",
2292 => x"0c873d0d",
2293 => x"0480e180",
2294 => x"08567580",
2295 => x"2ef03877",
2296 => x"76710c54",
2297 => x"74b00c87",
2298 => x"3d0d04fb",
2299 => x"3d0d800b",
2300 => x"80e1800c",
2301 => x"7a537952",
2302 => x"78518299",
2303 => x"3fb00855",
2304 => x"b008ff2e",
2305 => x"883874b0",
2306 => x"0c873d0d",
2307 => x"0480e180",
2308 => x"08567580",
2309 => x"2ef03877",
2310 => x"76710c54",
2311 => x"74b00c87",
2312 => x"3d0d04fe",
2313 => x"3d0d80e0",
2314 => x"f4085170",
2315 => x"8a3880e1",
2316 => x"847080e0",
2317 => x"f40c5170",
2318 => x"75125252",
2319 => x"ff537087",
2320 => x"fb808026",
2321 => x"88387080",
2322 => x"e0f40c71",
2323 => x"5372b00c",
2324 => x"843d0d04",
2325 => x"fd3d0d80",
2326 => x"0b80d0f8",
2327 => x"08545472",
2328 => x"812e9c38",
2329 => x"7380e0f8",
2330 => x"0cc0fb3f",
2331 => x"ffbf913f",
2332 => x"80e0cc52",
2333 => x"8151c386",
2334 => x"3fb00851",
2335 => x"85c63f72",
2336 => x"80e0f80c",
2337 => x"c0e03fff",
2338 => x"bef63f80",
2339 => x"e0cc5281",
2340 => x"51c2eb3f",
2341 => x"b0085185",
2342 => x"ab3f00ff",
2343 => x"39f53d0d",
2344 => x"7e6080e0",
2345 => x"f808705b",
2346 => x"585b5b75",
2347 => x"80c53877",
2348 => x"7a25a238",
2349 => x"771b7033",
2350 => x"7081ff06",
2351 => x"58585975",
2352 => x"8a2e9938",
2353 => x"7681ff06",
2354 => x"51ffbff9",
2355 => x"3f811858",
2356 => x"797824e0",
2357 => x"3879b00c",
2358 => x"8d3d0d04",
2359 => x"8d51ffbf",
2360 => x"e43f7833",
2361 => x"7081ff06",
2362 => x"5257ffbf",
2363 => x"d83f8118",
2364 => x"58de3979",
2365 => x"557a547d",
2366 => x"5385528d",
2367 => x"3dfc0551",
2368 => x"ffbebf3f",
2369 => x"b0085684",
2370 => x"b43f7bb0",
2371 => x"080c75b0",
2372 => x"0c8d3d0d",
2373 => x"04f63d0d",
2374 => x"7d7f80e0",
2375 => x"f808705b",
2376 => x"585a5a75",
2377 => x"80c43877",
2378 => x"7925b638",
2379 => x"ffbef13f",
2380 => x"b00881ff",
2381 => x"06708d32",
2382 => x"7030709f",
2383 => x"2a515157",
2384 => x"57768a2e",
2385 => x"80c63875",
2386 => x"802e80c0",
2387 => x"38771a56",
2388 => x"76763476",
2389 => x"51ffbeed",
2390 => x"3f811858",
2391 => x"787824cc",
2392 => x"38775675",
2393 => x"b00c8c3d",
2394 => x"0d047855",
2395 => x"79547c53",
2396 => x"84528c3d",
2397 => x"fc0551ff",
2398 => x"bdc83fb0",
2399 => x"085683bd",
2400 => x"3f7ab008",
2401 => x"0c75b00c",
2402 => x"8c3d0d04",
2403 => x"771a568a",
2404 => x"76348118",
2405 => x"588d51ff",
2406 => x"beab3f8a",
2407 => x"51ffbea5",
2408 => x"3f7756ff",
2409 => x"be39fb3d",
2410 => x"0d80e0f8",
2411 => x"08705654",
2412 => x"73883874",
2413 => x"b00c873d",
2414 => x"0d047753",
2415 => x"8352873d",
2416 => x"fc0551ff",
2417 => x"bcfc3fb0",
2418 => x"085482f1",
2419 => x"3f75b008",
2420 => x"0c73b00c",
2421 => x"873d0d04",
2422 => x"fa3d0d80",
2423 => x"e0f80880",
2424 => x"2ea3387a",
2425 => x"55795478",
2426 => x"53865288",
2427 => x"3dfc0551",
2428 => x"ffbccf3f",
2429 => x"b0085682",
2430 => x"c43f76b0",
2431 => x"080c75b0",
2432 => x"0c883d0d",
2433 => x"0482b63f",
2434 => x"9d0bb008",
2435 => x"0cff0bb0",
2436 => x"0c883d0d",
2437 => x"04fb3d0d",
2438 => x"77795656",
2439 => x"80705454",
2440 => x"7375259f",
2441 => x"38741010",
2442 => x"10f80552",
2443 => x"72167033",
2444 => x"70742b76",
2445 => x"078116f8",
2446 => x"16565656",
2447 => x"51517473",
2448 => x"24ea3873",
2449 => x"b00c873d",
2450 => x"0d04fc3d",
2451 => x"0d767855",
2452 => x"55bc5380",
2453 => x"527351f5",
2454 => x"be3f8452",
2455 => x"7451ffb5",
2456 => x"3fb00874",
2457 => x"23845284",
2458 => x"1551ffa9",
2459 => x"3fb00882",
2460 => x"15238452",
2461 => x"881551ff",
2462 => x"9c3fb008",
2463 => x"84150c84",
2464 => x"528c1551",
2465 => x"ff8f3fb0",
2466 => x"08881523",
2467 => x"84529015",
2468 => x"51ff823f",
2469 => x"b0088a15",
2470 => x"23845294",
2471 => x"1551fef5",
2472 => x"3fb0088c",
2473 => x"15238452",
2474 => x"981551fe",
2475 => x"e83fb008",
2476 => x"8e152388",
2477 => x"529c1551",
2478 => x"fedb3fb0",
2479 => x"0890150c",
2480 => x"863d0d04",
2481 => x"e93d0d6a",
2482 => x"80e0f808",
2483 => x"57577593",
2484 => x"3880c080",
2485 => x"0b84180c",
2486 => x"75ac180c",
2487 => x"75b00c99",
2488 => x"3d0d0489",
2489 => x"3d70556a",
2490 => x"54558a52",
2491 => x"993dffbc",
2492 => x"0551ffba",
2493 => x"cd3fb008",
2494 => x"77537552",
2495 => x"56fecb3f",
2496 => x"bc3f77b0",
2497 => x"080c75b0",
2498 => x"0c993d0d",
2499 => x"04fc3d0d",
2500 => x"815480e0",
2501 => x"f8088838",
2502 => x"73b00c86",
2503 => x"3d0d0476",
2504 => x"5397b952",
2505 => x"863dfc05",
2506 => x"51ffba96",
2507 => x"3fb00854",
2508 => x"8c3f74b0",
2509 => x"080c73b0",
2510 => x"0c863d0d",
2511 => x"0480d188",
2512 => x"08b00c04",
2513 => x"f73d0d7b",
2514 => x"80d18808",
2515 => x"82c81108",
2516 => x"5a545a77",
2517 => x"802e80da",
2518 => x"38818818",
2519 => x"841908ff",
2520 => x"0581712b",
2521 => x"59555980",
2522 => x"742480ea",
2523 => x"38807424",
2524 => x"b5387382",
2525 => x"2b781188",
2526 => x"05565681",
2527 => x"80190877",
2528 => x"06537280",
2529 => x"2eb63878",
2530 => x"16700853",
2531 => x"53795174",
2532 => x"0853722d",
2533 => x"ff14fc17",
2534 => x"fc177981",
2535 => x"2c5a5757",
2536 => x"54738025",
2537 => x"d6387708",
2538 => x"5877ffad",
2539 => x"3880d188",
2540 => x"0853bc13",
2541 => x"08a53879",
2542 => x"51f9df3f",
2543 => x"74085372",
2544 => x"2dff14fc",
2545 => x"17fc1779",
2546 => x"812c5a57",
2547 => x"57547380",
2548 => x"25ffa838",
2549 => x"d1398057",
2550 => x"ff933972",
2551 => x"51bc1308",
2552 => x"53722d79",
2553 => x"51f9b33f",
2554 => x"ff3d0d80",
2555 => x"e0d40bfc",
2556 => x"05700852",
2557 => x"5270ff2e",
2558 => x"9138702d",
2559 => x"fc127008",
2560 => x"525270ff",
2561 => x"2e098106",
2562 => x"f138833d",
2563 => x"0d0404ff",
2564 => x"babf3f04",
2565 => x"00ffffff",
2566 => x"ff00ffff",
2567 => x"ffff00ff",
2568 => x"ffffff00",
2569 => x"00000040",
2570 => x"30313233",
2571 => x"34353637",
2572 => x"38396162",
2573 => x"63646566",
2574 => x"00000000",
2575 => x"476f7420",
2576 => x"696e7465",
2577 => x"72727570",
2578 => x"740a0000",
2579 => x"633a0000",
2580 => x"733a0000",
2581 => x"4e6f2069",
2582 => x"6e746572",
2583 => x"72757074",
2584 => x"0a000000",
2585 => x"43000000",
2586 => x"64756d6d",
2587 => x"792e6578",
2588 => x"65000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"0000305c",
2593 => x"00002828",
2594 => x"0000288c",
2595 => x"00000000",
2596 => x"00002af4",
2597 => x"00002b50",
2598 => x"00002bac",
2599 => x"00000000",
2600 => x"00000000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00002864",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000001",
2638 => x"330eabcd",
2639 => x"1234e66d",
2640 => x"deec0005",
2641 => x"000b0000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000000",
2827 => x"00000000",
2828 => x"00000000",
2829 => x"00000000",
2830 => x"ffffffff",
2831 => x"00000000",
2832 => x"00020000",
2833 => x"00000000",
2834 => x"00000000",
2835 => x"00002c44",
2836 => x"00002c44",
2837 => x"00002c4c",
2838 => x"00002c4c",
2839 => x"00002c54",
2840 => x"00002c54",
2841 => x"00002c5c",
2842 => x"00002c5c",
2843 => x"00002c64",
2844 => x"00002c64",
2845 => x"00002c6c",
2846 => x"00002c6c",
2847 => x"00002c74",
2848 => x"00002c74",
2849 => x"00002c7c",
2850 => x"00002c7c",
2851 => x"00002c84",
2852 => x"00002c84",
2853 => x"00002c8c",
2854 => x"00002c8c",
2855 => x"00002c94",
2856 => x"00002c94",
2857 => x"00002c9c",
2858 => x"00002c9c",
2859 => x"00002ca4",
2860 => x"00002ca4",
2861 => x"00002cac",
2862 => x"00002cac",
2863 => x"00002cb4",
2864 => x"00002cb4",
2865 => x"00002cbc",
2866 => x"00002cbc",
2867 => x"00002cc4",
2868 => x"00002cc4",
2869 => x"00002ccc",
2870 => x"00002ccc",
2871 => x"00002cd4",
2872 => x"00002cd4",
2873 => x"00002cdc",
2874 => x"00002cdc",
2875 => x"00002ce4",
2876 => x"00002ce4",
2877 => x"00002cec",
2878 => x"00002cec",
2879 => x"00002cf4",
2880 => x"00002cf4",
2881 => x"00002cfc",
2882 => x"00002cfc",
2883 => x"00002d04",
2884 => x"00002d04",
2885 => x"00002d0c",
2886 => x"00002d0c",
2887 => x"00002d14",
2888 => x"00002d14",
2889 => x"00002d1c",
2890 => x"00002d1c",
2891 => x"00002d24",
2892 => x"00002d24",
2893 => x"00002d2c",
2894 => x"00002d2c",
2895 => x"00002d34",
2896 => x"00002d34",
2897 => x"00002d3c",
2898 => x"00002d3c",
2899 => x"00002d44",
2900 => x"00002d44",
2901 => x"00002d4c",
2902 => x"00002d4c",
2903 => x"00002d54",
2904 => x"00002d54",
2905 => x"00002d5c",
2906 => x"00002d5c",
2907 => x"00002d64",
2908 => x"00002d64",
2909 => x"00002d6c",
2910 => x"00002d6c",
2911 => x"00002d74",
2912 => x"00002d74",
2913 => x"00002d7c",
2914 => x"00002d7c",
2915 => x"00002d84",
2916 => x"00002d84",
2917 => x"00002d8c",
2918 => x"00002d8c",
2919 => x"00002d94",
2920 => x"00002d94",
2921 => x"00002d9c",
2922 => x"00002d9c",
2923 => x"00002da4",
2924 => x"00002da4",
2925 => x"00002dac",
2926 => x"00002dac",
2927 => x"00002db4",
2928 => x"00002db4",
2929 => x"00002dbc",
2930 => x"00002dbc",
2931 => x"00002dc4",
2932 => x"00002dc4",
2933 => x"00002dcc",
2934 => x"00002dcc",
2935 => x"00002dd4",
2936 => x"00002dd4",
2937 => x"00002ddc",
2938 => x"00002ddc",
2939 => x"00002de4",
2940 => x"00002de4",
2941 => x"00002dec",
2942 => x"00002dec",
2943 => x"00002df4",
2944 => x"00002df4",
2945 => x"00002dfc",
2946 => x"00002dfc",
2947 => x"00002e04",
2948 => x"00002e04",
2949 => x"00002e0c",
2950 => x"00002e0c",
2951 => x"00002e14",
2952 => x"00002e14",
2953 => x"00002e1c",
2954 => x"00002e1c",
2955 => x"00002e24",
2956 => x"00002e24",
2957 => x"00002e2c",
2958 => x"00002e2c",
2959 => x"00002e34",
2960 => x"00002e34",
2961 => x"00002e3c",
2962 => x"00002e3c",
2963 => x"00002e44",
2964 => x"00002e44",
2965 => x"00002e4c",
2966 => x"00002e4c",
2967 => x"00002e54",
2968 => x"00002e54",
2969 => x"00002e5c",
2970 => x"00002e5c",
2971 => x"00002e64",
2972 => x"00002e64",
2973 => x"00002e6c",
2974 => x"00002e6c",
2975 => x"00002e74",
2976 => x"00002e74",
2977 => x"00002e7c",
2978 => x"00002e7c",
2979 => x"00002e84",
2980 => x"00002e84",
2981 => x"00002e8c",
2982 => x"00002e8c",
2983 => x"00002e94",
2984 => x"00002e94",
2985 => x"00002e9c",
2986 => x"00002e9c",
2987 => x"00002ea4",
2988 => x"00002ea4",
2989 => x"00002eac",
2990 => x"00002eac",
2991 => x"00002eb4",
2992 => x"00002eb4",
2993 => x"00002ebc",
2994 => x"00002ebc",
2995 => x"00002ec4",
2996 => x"00002ec4",
2997 => x"00002ecc",
2998 => x"00002ecc",
2999 => x"00002ed4",
3000 => x"00002ed4",
3001 => x"00002edc",
3002 => x"00002edc",
3003 => x"00002ee4",
3004 => x"00002ee4",
3005 => x"00002eec",
3006 => x"00002eec",
3007 => x"00002ef4",
3008 => x"00002ef4",
3009 => x"00002efc",
3010 => x"00002efc",
3011 => x"00002f04",
3012 => x"00002f04",
3013 => x"00002f0c",
3014 => x"00002f0c",
3015 => x"00002f14",
3016 => x"00002f14",
3017 => x"00002f1c",
3018 => x"00002f1c",
3019 => x"00002f24",
3020 => x"00002f24",
3021 => x"00002f2c",
3022 => x"00002f2c",
3023 => x"00002f34",
3024 => x"00002f34",
3025 => x"00002f3c",
3026 => x"00002f3c",
3027 => x"00002f44",
3028 => x"00002f44",
3029 => x"00002f4c",
3030 => x"00002f4c",
3031 => x"00002f54",
3032 => x"00002f54",
3033 => x"00002f5c",
3034 => x"00002f5c",
3035 => x"00002f64",
3036 => x"00002f64",
3037 => x"00002f6c",
3038 => x"00002f6c",
3039 => x"00002f74",
3040 => x"00002f74",
3041 => x"00002f7c",
3042 => x"00002f7c",
3043 => x"00002f84",
3044 => x"00002f84",
3045 => x"00002f8c",
3046 => x"00002f8c",
3047 => x"00002f94",
3048 => x"00002f94",
3049 => x"00002f9c",
3050 => x"00002f9c",
3051 => x"00002fa4",
3052 => x"00002fa4",
3053 => x"00002fac",
3054 => x"00002fac",
3055 => x"00002fb4",
3056 => x"00002fb4",
3057 => x"00002fbc",
3058 => x"00002fbc",
3059 => x"00002fc4",
3060 => x"00002fc4",
3061 => x"00002fcc",
3062 => x"00002fcc",
3063 => x"00002fd4",
3064 => x"00002fd4",
3065 => x"00002fdc",
3066 => x"00002fdc",
3067 => x"00002fe4",
3068 => x"00002fe4",
3069 => x"00002fec",
3070 => x"00002fec",
3071 => x"00002ff4",
3072 => x"00002ff4",
3073 => x"00002ffc",
3074 => x"00002ffc",
3075 => x"00003004",
3076 => x"00003004",
3077 => x"0000300c",
3078 => x"0000300c",
3079 => x"00003014",
3080 => x"00003014",
3081 => x"0000301c",
3082 => x"0000301c",
3083 => x"00003024",
3084 => x"00003024",
3085 => x"0000302c",
3086 => x"0000302c",
3087 => x"00003034",
3088 => x"00003034",
3089 => x"0000303c",
3090 => x"0000303c",
3091 => x"00002868",
3092 => x"ffffffff",
3093 => x"00000000",
3094 => x"ffffffff",
3095 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

