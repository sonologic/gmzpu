------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cfe40c",
3 => x"3a0b0b80",
4 => x"c7ba0400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80ce",
162 => x"f4738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cfe00c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c6c03f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8ee82d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8db62d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80dfd0",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80df",
307 => x"d0085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480cf",
314 => x"e008802e",
315 => x"a43880cf",
316 => x"e408822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80dfd00c",
320 => x"82a0800b",
321 => x"80dfd40c",
322 => x"8290800b",
323 => x"80dfd80c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80dfd0",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"dfd40cf8",
330 => x"80808480",
331 => x"0b80dfd8",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80df",
335 => x"d00c80c0",
336 => x"a880940b",
337 => x"80dfd40c",
338 => x"80cf840b",
339 => x"80dfd80c",
340 => x"04ff3d0d",
341 => x"80dfdc33",
342 => x"5170a738",
343 => x"80cfec08",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"cfec0c70",
348 => x"2d80cfec",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80df",
352 => x"dc34833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80dfcc08",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"dfcc510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404803d",
366 => x"0d80dfe8",
367 => x"08811180",
368 => x"dfe80c51",
369 => x"800b8e80",
370 => x"800c823d",
371 => x"0d04f73d",
372 => x"0d7b5487",
373 => x"0b893d80",
374 => x"cff00858",
375 => x"58557417",
376 => x"748f0617",
377 => x"53537133",
378 => x"73347384",
379 => x"2aff1656",
380 => x"54748025",
381 => x"e938800b",
382 => x"8b3d3476",
383 => x"51878e3f",
384 => x"8b3d0d04",
385 => x"f33d0d80",
386 => x"cf9c5187",
387 => x"803f800b",
388 => x"8c80800c",
389 => x"8c808008",
390 => x"8c808408",
391 => x"80cfa053",
392 => x"595286e9",
393 => x"3f715487",
394 => x"0b8d3d80",
395 => x"cff00858",
396 => x"58557417",
397 => x"748f0617",
398 => x"53537133",
399 => x"73347384",
400 => x"2aff1656",
401 => x"54748025",
402 => x"e938800b",
403 => x"8f3d3476",
404 => x"5186ba3f",
405 => x"80cfa851",
406 => x"86b33f77",
407 => x"54870b80",
408 => x"cff0088b",
409 => x"3d595755",
410 => x"7417748f",
411 => x"06175458",
412 => x"72337834",
413 => x"73842aff",
414 => x"16565474",
415 => x"8025e938",
416 => x"800b8c3d",
417 => x"34765186",
418 => x"843f810b",
419 => x"8e80840c",
420 => x"80dfe808",
421 => x"5380dfe8",
422 => x"08547274",
423 => x"2e8f3880",
424 => x"cfb05185",
425 => x"e83f80df",
426 => x"e80853e9",
427 => x"3980cfc0",
428 => x"5185da3f",
429 => x"e039bc08",
430 => x"02bc0cf9",
431 => x"3d0d800b",
432 => x"bc08fc05",
433 => x"0cbc0888",
434 => x"05088025",
435 => x"ab38bc08",
436 => x"88050830",
437 => x"bc088805",
438 => x"0c800bbc",
439 => x"08f4050c",
440 => x"bc08fc05",
441 => x"08883881",
442 => x"0bbc08f4",
443 => x"050cbc08",
444 => x"f40508bc",
445 => x"08fc050c",
446 => x"bc088c05",
447 => x"088025ab",
448 => x"38bc088c",
449 => x"050830bc",
450 => x"088c050c",
451 => x"800bbc08",
452 => x"f0050cbc",
453 => x"08fc0508",
454 => x"8838810b",
455 => x"bc08f005",
456 => x"0cbc08f0",
457 => x"0508bc08",
458 => x"fc050c80",
459 => x"53bc088c",
460 => x"050852bc",
461 => x"08880508",
462 => x"5181a73f",
463 => x"b00870bc",
464 => x"08f8050c",
465 => x"54bc08fc",
466 => x"0508802e",
467 => x"8c38bc08",
468 => x"f8050830",
469 => x"bc08f805",
470 => x"0cbc08f8",
471 => x"050870b0",
472 => x"0c54893d",
473 => x"0dbc0c04",
474 => x"bc0802bc",
475 => x"0cfb3d0d",
476 => x"800bbc08",
477 => x"fc050cbc",
478 => x"08880508",
479 => x"80259338",
480 => x"bc088805",
481 => x"0830bc08",
482 => x"88050c81",
483 => x"0bbc08fc",
484 => x"050cbc08",
485 => x"8c050880",
486 => x"258c38bc",
487 => x"088c0508",
488 => x"30bc088c",
489 => x"050c8153",
490 => x"bc088c05",
491 => x"0852bc08",
492 => x"88050851",
493 => x"ad3fb008",
494 => x"70bc08f8",
495 => x"050c54bc",
496 => x"08fc0508",
497 => x"802e8c38",
498 => x"bc08f805",
499 => x"0830bc08",
500 => x"f8050cbc",
501 => x"08f80508",
502 => x"70b00c54",
503 => x"873d0dbc",
504 => x"0c04bc08",
505 => x"02bc0cfd",
506 => x"3d0d810b",
507 => x"bc08fc05",
508 => x"0c800bbc",
509 => x"08f8050c",
510 => x"bc088c05",
511 => x"08bc0888",
512 => x"050827ac",
513 => x"38bc08fc",
514 => x"0508802e",
515 => x"a338800b",
516 => x"bc088c05",
517 => x"08249938",
518 => x"bc088c05",
519 => x"0810bc08",
520 => x"8c050cbc",
521 => x"08fc0508",
522 => x"10bc08fc",
523 => x"050cc939",
524 => x"bc08fc05",
525 => x"08802e80",
526 => x"c938bc08",
527 => x"8c0508bc",
528 => x"08880508",
529 => x"26a138bc",
530 => x"08880508",
531 => x"bc088c05",
532 => x"0831bc08",
533 => x"88050cbc",
534 => x"08f80508",
535 => x"bc08fc05",
536 => x"0807bc08",
537 => x"f8050cbc",
538 => x"08fc0508",
539 => x"812abc08",
540 => x"fc050cbc",
541 => x"088c0508",
542 => x"812abc08",
543 => x"8c050cff",
544 => x"af39bc08",
545 => x"90050880",
546 => x"2e8f38bc",
547 => x"08880508",
548 => x"70bc08f4",
549 => x"050c518d",
550 => x"39bc08f8",
551 => x"050870bc",
552 => x"08f4050c",
553 => x"51bc08f4",
554 => x"0508b00c",
555 => x"853d0dbc",
556 => x"0c04fc3d",
557 => x"0d767079",
558 => x"7b555555",
559 => x"558f7227",
560 => x"8c387275",
561 => x"07830651",
562 => x"70802ea7",
563 => x"38ff1252",
564 => x"71ff2e98",
565 => x"38727081",
566 => x"05543374",
567 => x"70810556",
568 => x"34ff1252",
569 => x"71ff2e09",
570 => x"8106ea38",
571 => x"74b00c86",
572 => x"3d0d0474",
573 => x"51727084",
574 => x"05540871",
575 => x"70840553",
576 => x"0c727084",
577 => x"05540871",
578 => x"70840553",
579 => x"0c727084",
580 => x"05540871",
581 => x"70840553",
582 => x"0c727084",
583 => x"05540871",
584 => x"70840553",
585 => x"0cf01252",
586 => x"718f26c9",
587 => x"38837227",
588 => x"95387270",
589 => x"84055408",
590 => x"71708405",
591 => x"530cfc12",
592 => x"52718326",
593 => x"ed387054",
594 => x"ff8339f7",
595 => x"3d0d7c70",
596 => x"525380ca",
597 => x"3f7254b0",
598 => x"08550b0b",
599 => x"80cfcc56",
600 => x"8157b008",
601 => x"81055a8b",
602 => x"3de41159",
603 => x"538259f4",
604 => x"13527b88",
605 => x"11085253",
606 => x"81833fb0",
607 => x"083070b0",
608 => x"08079f2c",
609 => x"8a07b00c",
610 => x"538b3d0d",
611 => x"04ff3d0d",
612 => x"735280cf",
613 => x"f40851ff",
614 => x"b23f833d",
615 => x"0d04fd3d",
616 => x"0d757071",
617 => x"83065355",
618 => x"5270b838",
619 => x"71700870",
620 => x"09f7fbfd",
621 => x"ff120670",
622 => x"f8848281",
623 => x"80065151",
624 => x"5253709d",
625 => x"38841370",
626 => x"087009f7",
627 => x"fbfdff12",
628 => x"0670f884",
629 => x"82818006",
630 => x"51515253",
631 => x"70802ee5",
632 => x"38725271",
633 => x"33517080",
634 => x"2e8a3881",
635 => x"12703352",
636 => x"5270f838",
637 => x"717431b0",
638 => x"0c853d0d",
639 => x"04f23d0d",
640 => x"60628811",
641 => x"08705757",
642 => x"5f5a7480",
643 => x"2e818f38",
644 => x"8c1a2270",
645 => x"832a8132",
646 => x"70810651",
647 => x"55587386",
648 => x"38901a08",
649 => x"91387951",
650 => x"90a13fff",
651 => x"54b00880",
652 => x"ed388c1a",
653 => x"22587d08",
654 => x"57807883",
655 => x"ffff0670",
656 => x"812a7081",
657 => x"06515657",
658 => x"5573752e",
659 => x"80d73874",
660 => x"90387608",
661 => x"84180888",
662 => x"19595659",
663 => x"74802ef2",
664 => x"38745488",
665 => x"80752784",
666 => x"38888054",
667 => x"73537852",
668 => x"9c1a0851",
669 => x"a41a0854",
670 => x"732d800b",
671 => x"b0082582",
672 => x"e638b008",
673 => x"1975b008",
674 => x"317f8805",
675 => x"08b00831",
676 => x"70618805",
677 => x"0c565659",
678 => x"73ffb438",
679 => x"805473b0",
680 => x"0c903d0d",
681 => x"04758132",
682 => x"70810676",
683 => x"41515473",
684 => x"802e81c1",
685 => x"38749038",
686 => x"76088418",
687 => x"08881959",
688 => x"56597480",
689 => x"2ef23888",
690 => x"1a087883",
691 => x"ffff0670",
692 => x"892a7081",
693 => x"06515659",
694 => x"5673802e",
695 => x"82fa3875",
696 => x"75278d38",
697 => x"77872a70",
698 => x"81065154",
699 => x"7382b538",
700 => x"74762783",
701 => x"38745675",
702 => x"53785279",
703 => x"08518582",
704 => x"3f881a08",
705 => x"7631881b",
706 => x"0c790816",
707 => x"7a0c7456",
708 => x"75197577",
709 => x"317f8805",
710 => x"08783170",
711 => x"6188050c",
712 => x"56565973",
713 => x"802efef4",
714 => x"388c1a22",
715 => x"58ff8639",
716 => x"77785479",
717 => x"537b5256",
718 => x"84c83f88",
719 => x"1a087831",
720 => x"881b0c79",
721 => x"08187a0c",
722 => x"7c76315d",
723 => x"7c8e3879",
724 => x"518fdb3f",
725 => x"b008818f",
726 => x"38b0085f",
727 => x"75197577",
728 => x"317f8805",
729 => x"08783170",
730 => x"6188050c",
731 => x"56565973",
732 => x"802efea8",
733 => x"38748183",
734 => x"38760884",
735 => x"18088819",
736 => x"59565974",
737 => x"802ef238",
738 => x"74538a52",
739 => x"785182d3",
740 => x"3fb00879",
741 => x"3181055d",
742 => x"b0088438",
743 => x"81155d81",
744 => x"5f7c5874",
745 => x"7d278338",
746 => x"7458941a",
747 => x"08881b08",
748 => x"11575c80",
749 => x"7a085c54",
750 => x"901a087b",
751 => x"27833881",
752 => x"54757825",
753 => x"843873ba",
754 => x"387b7824",
755 => x"fee2387b",
756 => x"5378529c",
757 => x"1a0851a4",
758 => x"1a085473",
759 => x"2db00856",
760 => x"b0088024",
761 => x"fee2388c",
762 => x"1a2280c0",
763 => x"0754738c",
764 => x"1b23ff54",
765 => x"73b00c90",
766 => x"3d0d047e",
767 => x"ffa338ff",
768 => x"87397553",
769 => x"78527a51",
770 => x"82f83f79",
771 => x"08167a0c",
772 => x"79518e9a",
773 => x"3fb008cf",
774 => x"387c7631",
775 => x"5d7cfebc",
776 => x"38feac39",
777 => x"901a087a",
778 => x"08713176",
779 => x"1170565a",
780 => x"575280cf",
781 => x"f4085184",
782 => x"8c3fb008",
783 => x"802effa7",
784 => x"38b00890",
785 => x"1b0cb008",
786 => x"167a0c77",
787 => x"941b0c74",
788 => x"881b0c74",
789 => x"56fd9939",
790 => x"79085890",
791 => x"1a087827",
792 => x"83388154",
793 => x"75752784",
794 => x"3873b338",
795 => x"941a0856",
796 => x"75752680",
797 => x"d3387553",
798 => x"78529c1a",
799 => x"0851a41a",
800 => x"0854732d",
801 => x"b00856b0",
802 => x"088024fd",
803 => x"83388c1a",
804 => x"2280c007",
805 => x"54738c1b",
806 => x"23ff54fe",
807 => x"d7397553",
808 => x"78527751",
809 => x"81dc3f79",
810 => x"08167a0c",
811 => x"79518cfe",
812 => x"3fb00880",
813 => x"2efcd938",
814 => x"8c1a2280",
815 => x"c0075473",
816 => x"8c1b23ff",
817 => x"54fead39",
818 => x"74755479",
819 => x"53785256",
820 => x"81b03f88",
821 => x"1a087531",
822 => x"881b0c79",
823 => x"08157a0c",
824 => x"fcae39fa",
825 => x"3d0d7a79",
826 => x"028805a7",
827 => x"05335652",
828 => x"53837327",
829 => x"8a387083",
830 => x"06527180",
831 => x"2ea838ff",
832 => x"135372ff",
833 => x"2e973870",
834 => x"33527372",
835 => x"2e913881",
836 => x"11ff1454",
837 => x"5172ff2e",
838 => x"098106eb",
839 => x"38805170",
840 => x"b00c883d",
841 => x"0d047072",
842 => x"57558351",
843 => x"75828029",
844 => x"14ff1252",
845 => x"56708025",
846 => x"f3388373",
847 => x"27bf3874",
848 => x"08763270",
849 => x"09f7fbfd",
850 => x"ff120670",
851 => x"f8848281",
852 => x"80065151",
853 => x"5170802e",
854 => x"99387451",
855 => x"80527033",
856 => x"5773772e",
857 => x"ffb93881",
858 => x"11811353",
859 => x"51837227",
860 => x"ed38fc13",
861 => x"84165653",
862 => x"728326c3",
863 => x"387451fe",
864 => x"fe39fa3d",
865 => x"0d787a7c",
866 => x"72727257",
867 => x"57575956",
868 => x"56747627",
869 => x"b2387615",
870 => x"51757127",
871 => x"aa387077",
872 => x"17ff1454",
873 => x"555371ff",
874 => x"2e9638ff",
875 => x"14ff1454",
876 => x"54723374",
877 => x"34ff1252",
878 => x"71ff2e09",
879 => x"8106ec38",
880 => x"75b00c88",
881 => x"3d0d0476",
882 => x"8f269738",
883 => x"ff125271",
884 => x"ff2eed38",
885 => x"72708105",
886 => x"54337470",
887 => x"81055634",
888 => x"eb397476",
889 => x"07830651",
890 => x"70e23875",
891 => x"75545172",
892 => x"70840554",
893 => x"08717084",
894 => x"05530c72",
895 => x"70840554",
896 => x"08717084",
897 => x"05530c72",
898 => x"70840554",
899 => x"08717084",
900 => x"05530c72",
901 => x"70840554",
902 => x"08717084",
903 => x"05530cf0",
904 => x"1252718f",
905 => x"26c93883",
906 => x"72279538",
907 => x"72708405",
908 => x"54087170",
909 => x"8405530c",
910 => x"fc125271",
911 => x"8326ed38",
912 => x"7054ff88",
913 => x"39ef3d0d",
914 => x"63656740",
915 => x"5d427b80",
916 => x"2e84fa38",
917 => x"6151a5b4",
918 => x"3ff81c70",
919 => x"84120870",
920 => x"fc067062",
921 => x"8b0570f8",
922 => x"06415945",
923 => x"5b5c4157",
924 => x"96742782",
925 => x"c338807b",
926 => x"247e7c26",
927 => x"07598054",
928 => x"78742e09",
929 => x"810682a9",
930 => x"38777b25",
931 => x"81fc3877",
932 => x"1780d7b0",
933 => x"0b880508",
934 => x"5e567c76",
935 => x"2e84bd38",
936 => x"84160870",
937 => x"fe061784",
938 => x"11088106",
939 => x"51555573",
940 => x"828b3874",
941 => x"fc06597c",
942 => x"762e84dd",
943 => x"3877195f",
944 => x"7e7b2581",
945 => x"fd387981",
946 => x"06547382",
947 => x"bf387677",
948 => x"08318411",
949 => x"08fc0656",
950 => x"5a75802e",
951 => x"91387c76",
952 => x"2e84ea38",
953 => x"74191859",
954 => x"787b2584",
955 => x"89387980",
956 => x"2e829938",
957 => x"7715567a",
958 => x"76248290",
959 => x"388c1a08",
960 => x"881b0871",
961 => x"8c120c88",
962 => x"120c5579",
963 => x"76595788",
964 => x"1761fc05",
965 => x"575975a4",
966 => x"2685ef38",
967 => x"7b795555",
968 => x"93762780",
969 => x"c9387b70",
970 => x"84055d08",
971 => x"7c56790c",
972 => x"74708405",
973 => x"56088c18",
974 => x"0c901754",
975 => x"9b7627ae",
976 => x"38747084",
977 => x"05560874",
978 => x"0c747084",
979 => x"05560894",
980 => x"180c9817",
981 => x"54a37627",
982 => x"95387470",
983 => x"84055608",
984 => x"740c7470",
985 => x"84055608",
986 => x"9c180ca0",
987 => x"17547470",
988 => x"84055608",
989 => x"74708405",
990 => x"560c7470",
991 => x"84055608",
992 => x"74708405",
993 => x"560c7408",
994 => x"740c777b",
995 => x"3156758f",
996 => x"2680c938",
997 => x"84170881",
998 => x"06780784",
999 => x"180c7717",
1000 => x"84110881",
1001 => x"0784120c",
1002 => x"546151a2",
1003 => x"e03f8817",
1004 => x"5473b00c",
1005 => x"933d0d04",
1006 => x"905bfdba",
1007 => x"397856fe",
1008 => x"85398c16",
1009 => x"08881708",
1010 => x"718c120c",
1011 => x"88120c55",
1012 => x"7e707c31",
1013 => x"57588f76",
1014 => x"27ffb938",
1015 => x"7a178418",
1016 => x"0881067c",
1017 => x"0784190c",
1018 => x"76810784",
1019 => x"120c7611",
1020 => x"84110881",
1021 => x"0784120c",
1022 => x"55880552",
1023 => x"61518cf6",
1024 => x"3f6151a2",
1025 => x"883f8817",
1026 => x"54ffa639",
1027 => x"7d526151",
1028 => x"94f53fb0",
1029 => x"0859b008",
1030 => x"802e81a3",
1031 => x"38b008f8",
1032 => x"05608405",
1033 => x"08fe0661",
1034 => x"05555776",
1035 => x"742e83e6",
1036 => x"38fc1856",
1037 => x"75a42681",
1038 => x"aa387bb0",
1039 => x"08555593",
1040 => x"762780d8",
1041 => x"38747084",
1042 => x"055608b0",
1043 => x"08708405",
1044 => x"b00c0cb0",
1045 => x"08757084",
1046 => x"05570871",
1047 => x"70840553",
1048 => x"0c549b76",
1049 => x"27b63874",
1050 => x"70840556",
1051 => x"08747084",
1052 => x"05560c74",
1053 => x"70840556",
1054 => x"08747084",
1055 => x"05560ca3",
1056 => x"76279938",
1057 => x"74708405",
1058 => x"56087470",
1059 => x"8405560c",
1060 => x"74708405",
1061 => x"56087470",
1062 => x"8405560c",
1063 => x"74708405",
1064 => x"56087470",
1065 => x"8405560c",
1066 => x"74708405",
1067 => x"56087470",
1068 => x"8405560c",
1069 => x"7408740c",
1070 => x"7b526151",
1071 => x"8bb83f61",
1072 => x"51a0ca3f",
1073 => x"785473b0",
1074 => x"0c933d0d",
1075 => x"047d5261",
1076 => x"5193b43f",
1077 => x"b008b00c",
1078 => x"933d0d04",
1079 => x"84160855",
1080 => x"fbd13975",
1081 => x"537b52b0",
1082 => x"0851efc6",
1083 => x"3f7b5261",
1084 => x"518b833f",
1085 => x"ca398c16",
1086 => x"08881708",
1087 => x"718c120c",
1088 => x"88120c55",
1089 => x"8c1a0888",
1090 => x"1b08718c",
1091 => x"120c8812",
1092 => x"0c557979",
1093 => x"5957fbf7",
1094 => x"39771990",
1095 => x"1c555573",
1096 => x"7524fba2",
1097 => x"387a1770",
1098 => x"80d7b00b",
1099 => x"88050c75",
1100 => x"7c318107",
1101 => x"84120c5d",
1102 => x"84170881",
1103 => x"067b0784",
1104 => x"180c6151",
1105 => x"9fc73f88",
1106 => x"1754fce5",
1107 => x"39741918",
1108 => x"901c555d",
1109 => x"737d24fb",
1110 => x"95388c1a",
1111 => x"08881b08",
1112 => x"718c120c",
1113 => x"88120c55",
1114 => x"881a61fc",
1115 => x"05575975",
1116 => x"a42681ae",
1117 => x"387b7955",
1118 => x"55937627",
1119 => x"80c9387b",
1120 => x"7084055d",
1121 => x"087c5679",
1122 => x"0c747084",
1123 => x"0556088c",
1124 => x"1b0c901a",
1125 => x"549b7627",
1126 => x"ae387470",
1127 => x"84055608",
1128 => x"740c7470",
1129 => x"84055608",
1130 => x"941b0c98",
1131 => x"1a54a376",
1132 => x"27953874",
1133 => x"70840556",
1134 => x"08740c74",
1135 => x"70840556",
1136 => x"089c1b0c",
1137 => x"a01a5474",
1138 => x"70840556",
1139 => x"08747084",
1140 => x"05560c74",
1141 => x"70840556",
1142 => x"08747084",
1143 => x"05560c74",
1144 => x"08740c7a",
1145 => x"1a7080d7",
1146 => x"b00b8805",
1147 => x"0c7d7c31",
1148 => x"81078412",
1149 => x"0c54841a",
1150 => x"0881067b",
1151 => x"07841b0c",
1152 => x"61519e89",
1153 => x"3f7854fd",
1154 => x"bd397553",
1155 => x"7b527851",
1156 => x"eda03ffa",
1157 => x"f5398417",
1158 => x"08fc0618",
1159 => x"605858fa",
1160 => x"e9397553",
1161 => x"7b527851",
1162 => x"ed883f7a",
1163 => x"1a7080d7",
1164 => x"b00b8805",
1165 => x"0c7d7c31",
1166 => x"81078412",
1167 => x"0c54841a",
1168 => x"0881067b",
1169 => x"07841b0c",
1170 => x"ffb639fa",
1171 => x"3d0d7880",
1172 => x"cff40854",
1173 => x"55b81308",
1174 => x"802e81b5",
1175 => x"388c1522",
1176 => x"7083ffff",
1177 => x"0670832a",
1178 => x"81327081",
1179 => x"06515555",
1180 => x"5672802e",
1181 => x"80dc3873",
1182 => x"842a8132",
1183 => x"810657ff",
1184 => x"537680f6",
1185 => x"3873822a",
1186 => x"70810651",
1187 => x"5372802e",
1188 => x"b938b015",
1189 => x"08547380",
1190 => x"2e9c3880",
1191 => x"c0155373",
1192 => x"732e8f38",
1193 => x"735280cf",
1194 => x"f4085187",
1195 => x"c93f8c15",
1196 => x"225676b0",
1197 => x"160c75db",
1198 => x"0653728c",
1199 => x"1623800b",
1200 => x"84160c90",
1201 => x"1508750c",
1202 => x"72567588",
1203 => x"0753728c",
1204 => x"16239015",
1205 => x"08802e80",
1206 => x"c0388c15",
1207 => x"22708106",
1208 => x"5553739d",
1209 => x"3872812a",
1210 => x"70810651",
1211 => x"53728538",
1212 => x"94150854",
1213 => x"7388160c",
1214 => x"805372b0",
1215 => x"0c883d0d",
1216 => x"04800b88",
1217 => x"160c9415",
1218 => x"08309816",
1219 => x"0c8053ea",
1220 => x"39725182",
1221 => x"fb3ffec5",
1222 => x"3974518c",
1223 => x"e83f8c15",
1224 => x"22708106",
1225 => x"55537380",
1226 => x"2effba38",
1227 => x"d439f83d",
1228 => x"0d7a5877",
1229 => x"802e8199",
1230 => x"3880cff4",
1231 => x"0854b814",
1232 => x"08802e80",
1233 => x"ed388c18",
1234 => x"2270902b",
1235 => x"70902c70",
1236 => x"832a8132",
1237 => x"81065c51",
1238 => x"57547880",
1239 => x"cd389018",
1240 => x"08577680",
1241 => x"2e80c338",
1242 => x"77087731",
1243 => x"77790c76",
1244 => x"83067a58",
1245 => x"55557385",
1246 => x"38941808",
1247 => x"56758819",
1248 => x"0c807525",
1249 => x"a5387453",
1250 => x"76529c18",
1251 => x"0851a418",
1252 => x"0854732d",
1253 => x"800bb008",
1254 => x"2580c938",
1255 => x"b0081775",
1256 => x"b0083156",
1257 => x"57748024",
1258 => x"dd38800b",
1259 => x"b00c8a3d",
1260 => x"0d047351",
1261 => x"81da3f8c",
1262 => x"18227090",
1263 => x"2b70902c",
1264 => x"70832a81",
1265 => x"3281065c",
1266 => x"51575478",
1267 => x"dd38ff8e",
1268 => x"39a6ae52",
1269 => x"80cff408",
1270 => x"5189f13f",
1271 => x"b008b00c",
1272 => x"8a3d0d04",
1273 => x"8c182280",
1274 => x"c0075473",
1275 => x"8c1923ff",
1276 => x"0bb00c8a",
1277 => x"3d0d0480",
1278 => x"3d0d7251",
1279 => x"80710c80",
1280 => x"0b84120c",
1281 => x"800b8812",
1282 => x"0c028e05",
1283 => x"228c1223",
1284 => x"02920522",
1285 => x"8e122380",
1286 => x"0b90120c",
1287 => x"800b9412",
1288 => x"0c800b98",
1289 => x"120c709c",
1290 => x"120c80c2",
1291 => x"c20ba012",
1292 => x"0c80c38e",
1293 => x"0ba4120c",
1294 => x"80c48a0b",
1295 => x"a8120c80",
1296 => x"c4db0bac",
1297 => x"120c823d",
1298 => x"0d04fa3d",
1299 => x"0d797080",
1300 => x"dc298c11",
1301 => x"547a5356",
1302 => x"578cac3f",
1303 => x"b008b008",
1304 => x"5556b008",
1305 => x"802ea238",
1306 => x"b0088c05",
1307 => x"54800bb0",
1308 => x"080c76b0",
1309 => x"0884050c",
1310 => x"73b00888",
1311 => x"050c7453",
1312 => x"80527351",
1313 => x"97f73f75",
1314 => x"5473b00c",
1315 => x"883d0d04",
1316 => x"fc3d0d76",
1317 => x"aba30bbc",
1318 => x"120c5581",
1319 => x"0bb8160c",
1320 => x"800b84dc",
1321 => x"160c830b",
1322 => x"84e0160c",
1323 => x"84e81584",
1324 => x"e4160c74",
1325 => x"54805384",
1326 => x"52841508",
1327 => x"51feb83f",
1328 => x"74548153",
1329 => x"89528815",
1330 => x"0851feab",
1331 => x"3f745482",
1332 => x"538a528c",
1333 => x"150851fe",
1334 => x"9e3f863d",
1335 => x"0d04f93d",
1336 => x"0d7980cf",
1337 => x"f4085457",
1338 => x"b8130880",
1339 => x"2e80c838",
1340 => x"84dc1356",
1341 => x"88160884",
1342 => x"1708ff05",
1343 => x"55558074",
1344 => x"249f388c",
1345 => x"15227090",
1346 => x"2b70902c",
1347 => x"51545872",
1348 => x"802e80ca",
1349 => x"3880dc15",
1350 => x"ff155555",
1351 => x"738025e3",
1352 => x"38750853",
1353 => x"72802e9f",
1354 => x"38725688",
1355 => x"16088417",
1356 => x"08ff0555",
1357 => x"55c83972",
1358 => x"51fed53f",
1359 => x"80cff408",
1360 => x"84dc0556",
1361 => x"ffae3984",
1362 => x"527651fd",
1363 => x"fd3fb008",
1364 => x"760cb008",
1365 => x"802e80c0",
1366 => x"38b00856",
1367 => x"ce39810b",
1368 => x"8c162372",
1369 => x"750c7288",
1370 => x"160c7284",
1371 => x"160c7290",
1372 => x"160c7294",
1373 => x"160c7298",
1374 => x"160cff0b",
1375 => x"8e162372",
1376 => x"b0160c72",
1377 => x"b4160c72",
1378 => x"80c4160c",
1379 => x"7280c816",
1380 => x"0c74b00c",
1381 => x"893d0d04",
1382 => x"8c770c80",
1383 => x"0bb00c89",
1384 => x"3d0d04ff",
1385 => x"3d0da6ae",
1386 => x"52735186",
1387 => x"9f3f833d",
1388 => x"0d04803d",
1389 => x"0d80cff4",
1390 => x"0851e83f",
1391 => x"823d0d04",
1392 => x"fb3d0d77",
1393 => x"70525696",
1394 => x"c33f80d7",
1395 => x"b00b8805",
1396 => x"08841108",
1397 => x"fc06707b",
1398 => x"319fef05",
1399 => x"e08006e0",
1400 => x"80055656",
1401 => x"53a08074",
1402 => x"24943880",
1403 => x"52755196",
1404 => x"9d3f80d7",
1405 => x"b8081553",
1406 => x"72b0082e",
1407 => x"8f387551",
1408 => x"968b3f80",
1409 => x"5372b00c",
1410 => x"873d0d04",
1411 => x"73305275",
1412 => x"5195fb3f",
1413 => x"b008ff2e",
1414 => x"a83880d7",
1415 => x"b00b8805",
1416 => x"08757531",
1417 => x"81078412",
1418 => x"0c5380d6",
1419 => x"f4087431",
1420 => x"80d6f40c",
1421 => x"755195d5",
1422 => x"3f810bb0",
1423 => x"0c873d0d",
1424 => x"04805275",
1425 => x"5195c73f",
1426 => x"80d7b00b",
1427 => x"880508b0",
1428 => x"08713156",
1429 => x"538f7525",
1430 => x"ffa438b0",
1431 => x"0880d7a4",
1432 => x"083180d6",
1433 => x"f40c7481",
1434 => x"0784140c",
1435 => x"7551959d",
1436 => x"3f8053ff",
1437 => x"9039f63d",
1438 => x"0d7c7e54",
1439 => x"5b72802e",
1440 => x"8283387a",
1441 => x"5195853f",
1442 => x"f8138411",
1443 => x"0870fe06",
1444 => x"70138411",
1445 => x"08fc065d",
1446 => x"58595458",
1447 => x"80d7b808",
1448 => x"752e82de",
1449 => x"38788416",
1450 => x"0c807381",
1451 => x"06545a72",
1452 => x"7a2e81d5",
1453 => x"38781584",
1454 => x"11088106",
1455 => x"515372a0",
1456 => x"38781757",
1457 => x"7981e638",
1458 => x"88150853",
1459 => x"7280d7b8",
1460 => x"2e82f938",
1461 => x"8c150870",
1462 => x"8c150c73",
1463 => x"88120c56",
1464 => x"76810784",
1465 => x"190c7618",
1466 => x"77710c53",
1467 => x"79819138",
1468 => x"83ff7727",
1469 => x"81c83876",
1470 => x"892a7783",
1471 => x"2a565372",
1472 => x"802ebf38",
1473 => x"76862ab8",
1474 => x"05558473",
1475 => x"27b43880",
1476 => x"db135594",
1477 => x"7327ab38",
1478 => x"768c2a80",
1479 => x"ee055580",
1480 => x"d473279e",
1481 => x"38768f2a",
1482 => x"80f70555",
1483 => x"82d47327",
1484 => x"91387692",
1485 => x"2a80fc05",
1486 => x"558ad473",
1487 => x"27843880",
1488 => x"fe557410",
1489 => x"101080d7",
1490 => x"b0058811",
1491 => x"08555673",
1492 => x"762e82b3",
1493 => x"38841408",
1494 => x"fc065376",
1495 => x"73278d38",
1496 => x"88140854",
1497 => x"73762e09",
1498 => x"8106ea38",
1499 => x"8c140870",
1500 => x"8c1a0c74",
1501 => x"881a0c78",
1502 => x"88120c56",
1503 => x"778c150c",
1504 => x"7a519389",
1505 => x"3f8c3d0d",
1506 => x"04770878",
1507 => x"71315977",
1508 => x"05881908",
1509 => x"54577280",
1510 => x"d7b82e80",
1511 => x"e0388c18",
1512 => x"08708c15",
1513 => x"0c738812",
1514 => x"0c56fe89",
1515 => x"39881508",
1516 => x"8c160870",
1517 => x"8c130c57",
1518 => x"88170cfe",
1519 => x"a3397683",
1520 => x"2a705455",
1521 => x"80752481",
1522 => x"98387282",
1523 => x"2c81712b",
1524 => x"80d7b408",
1525 => x"0780d7b0",
1526 => x"0b84050c",
1527 => x"53741010",
1528 => x"1080d7b0",
1529 => x"05881108",
1530 => x"5556758c",
1531 => x"190c7388",
1532 => x"190c7788",
1533 => x"170c778c",
1534 => x"150cff84",
1535 => x"39815afd",
1536 => x"b4397817",
1537 => x"73810654",
1538 => x"57729838",
1539 => x"77087871",
1540 => x"31597705",
1541 => x"8c190888",
1542 => x"1a08718c",
1543 => x"120c8812",
1544 => x"0c575776",
1545 => x"81078419",
1546 => x"0c7780d7",
1547 => x"b00b8805",
1548 => x"0c80d7ac",
1549 => x"087726fe",
1550 => x"c73880d7",
1551 => x"a808527a",
1552 => x"51fafd3f",
1553 => x"7a5191c5",
1554 => x"3ffeba39",
1555 => x"81788c15",
1556 => x"0c788815",
1557 => x"0c738c1a",
1558 => x"0c73881a",
1559 => x"0c5afd80",
1560 => x"39831570",
1561 => x"822c8171",
1562 => x"2b80d7b4",
1563 => x"080780d7",
1564 => x"b00b8405",
1565 => x"0c515374",
1566 => x"10101080",
1567 => x"d7b00588",
1568 => x"11085556",
1569 => x"fee43974",
1570 => x"53807524",
1571 => x"a7387282",
1572 => x"2c81712b",
1573 => x"80d7b408",
1574 => x"0780d7b0",
1575 => x"0b84050c",
1576 => x"53758c19",
1577 => x"0c738819",
1578 => x"0c778817",
1579 => x"0c778c15",
1580 => x"0cfdcd39",
1581 => x"83157082",
1582 => x"2c81712b",
1583 => x"80d7b408",
1584 => x"0780d7b0",
1585 => x"0b84050c",
1586 => x"5153d639",
1587 => x"f93d0d79",
1588 => x"7b585380",
1589 => x"0b80cff4",
1590 => x"08535672",
1591 => x"722e80c0",
1592 => x"3884dc13",
1593 => x"5574762e",
1594 => x"b7388815",
1595 => x"08841608",
1596 => x"ff055454",
1597 => x"8073249d",
1598 => x"388c1422",
1599 => x"70902b70",
1600 => x"902c5153",
1601 => x"587180d8",
1602 => x"3880dc14",
1603 => x"ff145454",
1604 => x"728025e5",
1605 => x"38740855",
1606 => x"74d03880",
1607 => x"cff40852",
1608 => x"84dc1255",
1609 => x"74802eb1",
1610 => x"38881508",
1611 => x"841608ff",
1612 => x"05545480",
1613 => x"73249c38",
1614 => x"8c142270",
1615 => x"902b7090",
1616 => x"2c515358",
1617 => x"71ad3880",
1618 => x"dc14ff14",
1619 => x"54547280",
1620 => x"25e63874",
1621 => x"085574d1",
1622 => x"3875b00c",
1623 => x"893d0d04",
1624 => x"7351762d",
1625 => x"75b00807",
1626 => x"80dc15ff",
1627 => x"15555556",
1628 => x"ff9e3973",
1629 => x"51762d75",
1630 => x"b0080780",
1631 => x"dc15ff15",
1632 => x"555556ca",
1633 => x"39ea3d0d",
1634 => x"688c1122",
1635 => x"70812a81",
1636 => x"06575856",
1637 => x"7480e438",
1638 => x"8e162270",
1639 => x"902b7090",
1640 => x"2c515558",
1641 => x"807424b1",
1642 => x"38983dc4",
1643 => x"05537352",
1644 => x"80cff408",
1645 => x"5192ac3f",
1646 => x"800bb008",
1647 => x"24973879",
1648 => x"83e08006",
1649 => x"547380c0",
1650 => x"802e818f",
1651 => x"38738280",
1652 => x"802e8191",
1653 => x"388c1622",
1654 => x"57769080",
1655 => x"0754738c",
1656 => x"17238880",
1657 => x"5280cff4",
1658 => x"0851819b",
1659 => x"3fb0089d",
1660 => x"388c1622",
1661 => x"82075473",
1662 => x"8c172380",
1663 => x"c3167077",
1664 => x"0c90170c",
1665 => x"810b9417",
1666 => x"0c983d0d",
1667 => x"0480cff4",
1668 => x"08aba30b",
1669 => x"bc120c54",
1670 => x"8c162281",
1671 => x"80075473",
1672 => x"8c1723b0",
1673 => x"08760cb0",
1674 => x"0890170c",
1675 => x"88800b94",
1676 => x"170c7480",
1677 => x"2ed3388e",
1678 => x"16227090",
1679 => x"2b70902c",
1680 => x"53555898",
1681 => x"a63fb008",
1682 => x"802effbd",
1683 => x"388c1622",
1684 => x"81075473",
1685 => x"8c172398",
1686 => x"3d0d0481",
1687 => x"0b8c1722",
1688 => x"5855fef5",
1689 => x"39a81608",
1690 => x"80c48a2e",
1691 => x"098106fe",
1692 => x"e4388c16",
1693 => x"22888007",
1694 => x"54738c17",
1695 => x"2388800b",
1696 => x"80cc170c",
1697 => x"fedc39f3",
1698 => x"3d0d7f61",
1699 => x"8b1170f8",
1700 => x"065c5555",
1701 => x"5e729626",
1702 => x"83389059",
1703 => x"80792474",
1704 => x"7a260753",
1705 => x"80547274",
1706 => x"2e098106",
1707 => x"80cb387d",
1708 => x"518cd93f",
1709 => x"7883f726",
1710 => x"80c63878",
1711 => x"832a7010",
1712 => x"101080d7",
1713 => x"b0058c11",
1714 => x"0859595a",
1715 => x"76782e83",
1716 => x"b0388417",
1717 => x"08fc0656",
1718 => x"8c170888",
1719 => x"1808718c",
1720 => x"120c8812",
1721 => x"0c587517",
1722 => x"84110881",
1723 => x"0784120c",
1724 => x"537d518c",
1725 => x"983f8817",
1726 => x"5473b00c",
1727 => x"8f3d0d04",
1728 => x"78892a79",
1729 => x"832a5b53",
1730 => x"72802ebf",
1731 => x"3878862a",
1732 => x"b8055a84",
1733 => x"7327b438",
1734 => x"80db135a",
1735 => x"947327ab",
1736 => x"38788c2a",
1737 => x"80ee055a",
1738 => x"80d47327",
1739 => x"9e38788f",
1740 => x"2a80f705",
1741 => x"5a82d473",
1742 => x"27913878",
1743 => x"922a80fc",
1744 => x"055a8ad4",
1745 => x"73278438",
1746 => x"80fe5a79",
1747 => x"10101080",
1748 => x"d7b0058c",
1749 => x"11085855",
1750 => x"76752ea3",
1751 => x"38841708",
1752 => x"fc06707a",
1753 => x"31555673",
1754 => x"8f2488d5",
1755 => x"38738025",
1756 => x"fee6388c",
1757 => x"17085776",
1758 => x"752e0981",
1759 => x"06df3881",
1760 => x"1a5a80d7",
1761 => x"c0085776",
1762 => x"80d7b82e",
1763 => x"82c03884",
1764 => x"1708fc06",
1765 => x"707a3155",
1766 => x"56738f24",
1767 => x"81f93880",
1768 => x"d7b80b80",
1769 => x"d7c40c80",
1770 => x"d7b80b80",
1771 => x"d7c00c73",
1772 => x"8025feb2",
1773 => x"3883ff76",
1774 => x"2783df38",
1775 => x"75892a76",
1776 => x"832a5553",
1777 => x"72802ebf",
1778 => x"3875862a",
1779 => x"b8055484",
1780 => x"7327b438",
1781 => x"80db1354",
1782 => x"947327ab",
1783 => x"38758c2a",
1784 => x"80ee0554",
1785 => x"80d47327",
1786 => x"9e38758f",
1787 => x"2a80f705",
1788 => x"5482d473",
1789 => x"27913875",
1790 => x"922a80fc",
1791 => x"05548ad4",
1792 => x"73278438",
1793 => x"80fe5473",
1794 => x"10101080",
1795 => x"d7b00588",
1796 => x"11085658",
1797 => x"74782e86",
1798 => x"cf388415",
1799 => x"08fc0653",
1800 => x"7573278d",
1801 => x"38881508",
1802 => x"5574782e",
1803 => x"098106ea",
1804 => x"388c1508",
1805 => x"80d7b00b",
1806 => x"84050871",
1807 => x"8c1a0c76",
1808 => x"881a0c78",
1809 => x"88130c78",
1810 => x"8c180c5d",
1811 => x"58795380",
1812 => x"7a2483e6",
1813 => x"3872822c",
1814 => x"81712b5c",
1815 => x"537a7c26",
1816 => x"8198387b",
1817 => x"7b065372",
1818 => x"82f13879",
1819 => x"fc068405",
1820 => x"5a7a1070",
1821 => x"7d06545b",
1822 => x"7282e038",
1823 => x"841a5af1",
1824 => x"3988178c",
1825 => x"11085858",
1826 => x"76782e09",
1827 => x"8106fcc2",
1828 => x"38821a5a",
1829 => x"fdec3978",
1830 => x"17798107",
1831 => x"84190c70",
1832 => x"80d7c40c",
1833 => x"7080d7c0",
1834 => x"0c80d7b8",
1835 => x"0b8c120c",
1836 => x"8c110888",
1837 => x"120c7481",
1838 => x"0784120c",
1839 => x"74117571",
1840 => x"0c51537d",
1841 => x"5188c63f",
1842 => x"881754fc",
1843 => x"ac3980d7",
1844 => x"b00b8405",
1845 => x"087a545c",
1846 => x"798025fe",
1847 => x"f83882da",
1848 => x"397a097c",
1849 => x"067080d7",
1850 => x"b00b8405",
1851 => x"0c5c7a10",
1852 => x"5b7a7c26",
1853 => x"85387a85",
1854 => x"b83880d7",
1855 => x"b00b8805",
1856 => x"08708412",
1857 => x"08fc0670",
1858 => x"7c317c72",
1859 => x"268f7225",
1860 => x"0757575c",
1861 => x"5d557280",
1862 => x"2e80db38",
1863 => x"797a1680",
1864 => x"d7a8081b",
1865 => x"90115a55",
1866 => x"575b80d7",
1867 => x"a408ff2e",
1868 => x"8838a08f",
1869 => x"13e08006",
1870 => x"5776527d",
1871 => x"5187cf3f",
1872 => x"b00854b0",
1873 => x"08ff2e90",
1874 => x"38b00876",
1875 => x"27829938",
1876 => x"7480d7b0",
1877 => x"2e829138",
1878 => x"80d7b00b",
1879 => x"88050855",
1880 => x"841508fc",
1881 => x"06707a31",
1882 => x"7a72268f",
1883 => x"72250752",
1884 => x"55537283",
1885 => x"e6387479",
1886 => x"81078417",
1887 => x"0c791670",
1888 => x"80d7b00b",
1889 => x"88050c75",
1890 => x"81078412",
1891 => x"0c547e52",
1892 => x"5786fa3f",
1893 => x"881754fa",
1894 => x"e0397583",
1895 => x"2a705454",
1896 => x"80742481",
1897 => x"9b387282",
1898 => x"2c81712b",
1899 => x"80d7b408",
1900 => x"077080d7",
1901 => x"b00b8405",
1902 => x"0c751010",
1903 => x"1080d7b0",
1904 => x"05881108",
1905 => x"585a5d53",
1906 => x"778c180c",
1907 => x"7488180c",
1908 => x"7688190c",
1909 => x"768c160c",
1910 => x"fcf33979",
1911 => x"7a101010",
1912 => x"80d7b005",
1913 => x"7057595d",
1914 => x"8c150857",
1915 => x"76752ea3",
1916 => x"38841708",
1917 => x"fc06707a",
1918 => x"31555673",
1919 => x"8f2483ca",
1920 => x"38738025",
1921 => x"8481388c",
1922 => x"17085776",
1923 => x"752e0981",
1924 => x"06df3888",
1925 => x"15811b70",
1926 => x"8306555b",
1927 => x"5572c938",
1928 => x"7c830653",
1929 => x"72802efd",
1930 => x"b838ff1d",
1931 => x"f819595d",
1932 => x"88180878",
1933 => x"2eea38fd",
1934 => x"b539831a",
1935 => x"53fc9639",
1936 => x"83147082",
1937 => x"2c81712b",
1938 => x"80d7b408",
1939 => x"077080d7",
1940 => x"b00b8405",
1941 => x"0c761010",
1942 => x"1080d7b0",
1943 => x"05881108",
1944 => x"595b5e51",
1945 => x"53fee139",
1946 => x"80d6f408",
1947 => x"1758b008",
1948 => x"762e818d",
1949 => x"3880d7a4",
1950 => x"08ff2e83",
1951 => x"ec387376",
1952 => x"311880d6",
1953 => x"f40c7387",
1954 => x"06705753",
1955 => x"72802e88",
1956 => x"38887331",
1957 => x"70155556",
1958 => x"76149fff",
1959 => x"06a08071",
1960 => x"31177054",
1961 => x"7f535753",
1962 => x"84e43fb0",
1963 => x"0853b008",
1964 => x"ff2e81a0",
1965 => x"3880d6f4",
1966 => x"08167080",
1967 => x"d6f40c74",
1968 => x"7580d7b0",
1969 => x"0b88050c",
1970 => x"74763118",
1971 => x"70810751",
1972 => x"5556587b",
1973 => x"80d7b02e",
1974 => x"839c3879",
1975 => x"8f2682cb",
1976 => x"38810b84",
1977 => x"150c8415",
1978 => x"08fc0670",
1979 => x"7a317a72",
1980 => x"268f7225",
1981 => x"07525553",
1982 => x"72802efc",
1983 => x"f93880db",
1984 => x"39b0089f",
1985 => x"ff065372",
1986 => x"feeb3877",
1987 => x"80d6f40c",
1988 => x"80d7b00b",
1989 => x"8805087b",
1990 => x"18810784",
1991 => x"120c5580",
1992 => x"d7a00878",
1993 => x"27863877",
1994 => x"80d7a00c",
1995 => x"80d79c08",
1996 => x"7827fcac",
1997 => x"387780d7",
1998 => x"9c0c8415",
1999 => x"08fc0670",
2000 => x"7a317a72",
2001 => x"268f7225",
2002 => x"07525553",
2003 => x"72802efc",
2004 => x"a5388839",
2005 => x"80745456",
2006 => x"fedb397d",
2007 => x"5183ae3f",
2008 => x"800bb00c",
2009 => x"8f3d0d04",
2010 => x"73538074",
2011 => x"24a93872",
2012 => x"822c8171",
2013 => x"2b80d7b4",
2014 => x"08077080",
2015 => x"d7b00b84",
2016 => x"050c5d53",
2017 => x"778c180c",
2018 => x"7488180c",
2019 => x"7688190c",
2020 => x"768c160c",
2021 => x"f9b73983",
2022 => x"1470822c",
2023 => x"81712b80",
2024 => x"d7b40807",
2025 => x"7080d7b0",
2026 => x"0b84050c",
2027 => x"5e5153d4",
2028 => x"397b7b06",
2029 => x"5372fca3",
2030 => x"38841a7b",
2031 => x"105c5af1",
2032 => x"39ff1a81",
2033 => x"11515af7",
2034 => x"b9397817",
2035 => x"79810784",
2036 => x"190c8c18",
2037 => x"08881908",
2038 => x"718c120c",
2039 => x"88120c59",
2040 => x"7080d7c4",
2041 => x"0c7080d7",
2042 => x"c00c80d7",
2043 => x"b80b8c12",
2044 => x"0c8c1108",
2045 => x"88120c74",
2046 => x"81078412",
2047 => x"0c741175",
2048 => x"710c5153",
2049 => x"f9bd3975",
2050 => x"17841108",
2051 => x"81078412",
2052 => x"0c538c17",
2053 => x"08881808",
2054 => x"718c120c",
2055 => x"88120c58",
2056 => x"7d5181e9",
2057 => x"3f881754",
2058 => x"f5cf3972",
2059 => x"84150cf4",
2060 => x"1af80670",
2061 => x"841e0881",
2062 => x"0607841e",
2063 => x"0c701d54",
2064 => x"5b850b84",
2065 => x"140c850b",
2066 => x"88140c8f",
2067 => x"7b27fdcf",
2068 => x"38881c52",
2069 => x"7d51ec9e",
2070 => x"3f80d7b0",
2071 => x"0b880508",
2072 => x"80d6f408",
2073 => x"5955fdb7",
2074 => x"397780d6",
2075 => x"f40c7380",
2076 => x"d7a40cfc",
2077 => x"91397284",
2078 => x"150cfda3",
2079 => x"39fc3d0d",
2080 => x"76797102",
2081 => x"8c059f05",
2082 => x"33575553",
2083 => x"55837227",
2084 => x"8a387483",
2085 => x"06517080",
2086 => x"2ea238ff",
2087 => x"125271ff",
2088 => x"2e933873",
2089 => x"73708105",
2090 => x"5534ff12",
2091 => x"5271ff2e",
2092 => x"098106ef",
2093 => x"3874b00c",
2094 => x"863d0d04",
2095 => x"7474882b",
2096 => x"75077071",
2097 => x"902b0751",
2098 => x"54518f72",
2099 => x"27a53872",
2100 => x"71708405",
2101 => x"530c7271",
2102 => x"70840553",
2103 => x"0c727170",
2104 => x"8405530c",
2105 => x"72717084",
2106 => x"05530cf0",
2107 => x"1252718f",
2108 => x"26dd3883",
2109 => x"72279038",
2110 => x"72717084",
2111 => x"05530cfc",
2112 => x"12527183",
2113 => x"26f23870",
2114 => x"53ff9039",
2115 => x"0404fd3d",
2116 => x"0d800b80",
2117 => x"dfec0c76",
2118 => x"5184ee3f",
2119 => x"b00853b0",
2120 => x"08ff2e88",
2121 => x"3872b00c",
2122 => x"853d0d04",
2123 => x"80dfec08",
2124 => x"5473802e",
2125 => x"f0387574",
2126 => x"710c5272",
2127 => x"b00c853d",
2128 => x"0d04f93d",
2129 => x"0d797c55",
2130 => x"7b548e11",
2131 => x"2270902b",
2132 => x"70902c55",
2133 => x"5780cff4",
2134 => x"08535856",
2135 => x"83f33fb0",
2136 => x"0857800b",
2137 => x"b0082493",
2138 => x"3880d016",
2139 => x"08b00805",
2140 => x"80d0170c",
2141 => x"76b00c89",
2142 => x"3d0d048c",
2143 => x"162283df",
2144 => x"ff065574",
2145 => x"8c172376",
2146 => x"b00c893d",
2147 => x"0d04fa3d",
2148 => x"0d788c11",
2149 => x"2270882a",
2150 => x"70810651",
2151 => x"57585674",
2152 => x"a9388c16",
2153 => x"2283dfff",
2154 => x"0655748c",
2155 => x"17237a54",
2156 => x"79538e16",
2157 => x"2270902b",
2158 => x"70902c54",
2159 => x"5680cff4",
2160 => x"08525681",
2161 => x"b23f883d",
2162 => x"0d048254",
2163 => x"80538e16",
2164 => x"2270902b",
2165 => x"70902c54",
2166 => x"5680cff4",
2167 => x"08525782",
2168 => x"b83f8c16",
2169 => x"2283dfff",
2170 => x"0655748c",
2171 => x"17237a54",
2172 => x"79538e16",
2173 => x"2270902b",
2174 => x"70902c54",
2175 => x"5680cff4",
2176 => x"08525680",
2177 => x"f23f883d",
2178 => x"0d04f93d",
2179 => x"0d797c55",
2180 => x"7b548e11",
2181 => x"2270902b",
2182 => x"70902c55",
2183 => x"5780cff4",
2184 => x"08535856",
2185 => x"81f33fb0",
2186 => x"0857b008",
2187 => x"ff2e9938",
2188 => x"8c1622a0",
2189 => x"80075574",
2190 => x"8c1723b0",
2191 => x"0880d017",
2192 => x"0c76b00c",
2193 => x"893d0d04",
2194 => x"8c162283",
2195 => x"dfff0655",
2196 => x"748c1723",
2197 => x"76b00c89",
2198 => x"3d0d04fe",
2199 => x"3d0d748e",
2200 => x"11227090",
2201 => x"2b70902c",
2202 => x"55515153",
2203 => x"80cff408",
2204 => x"51bd3f84",
2205 => x"3d0d04fb",
2206 => x"3d0d800b",
2207 => x"80dfec0c",
2208 => x"7a537952",
2209 => x"785182f9",
2210 => x"3fb00855",
2211 => x"b008ff2e",
2212 => x"883874b0",
2213 => x"0c873d0d",
2214 => x"0480dfec",
2215 => x"08567580",
2216 => x"2ef03877",
2217 => x"76710c54",
2218 => x"74b00c87",
2219 => x"3d0d04fd",
2220 => x"3d0d800b",
2221 => x"80dfec0c",
2222 => x"765184c8",
2223 => x"3fb00853",
2224 => x"b008ff2e",
2225 => x"883872b0",
2226 => x"0c853d0d",
2227 => x"0480dfec",
2228 => x"08547380",
2229 => x"2ef03875",
2230 => x"74710c52",
2231 => x"72b00c85",
2232 => x"3d0d04fc",
2233 => x"3d0d800b",
2234 => x"80dfec0c",
2235 => x"78527751",
2236 => x"86b03fb0",
2237 => x"0854b008",
2238 => x"ff2e8838",
2239 => x"73b00c86",
2240 => x"3d0d0480",
2241 => x"dfec0855",
2242 => x"74802ef0",
2243 => x"38767571",
2244 => x"0c5373b0",
2245 => x"0c863d0d",
2246 => x"04fb3d0d",
2247 => x"800b80df",
2248 => x"ec0c7a53",
2249 => x"79527851",
2250 => x"848c3fb0",
2251 => x"0855b008",
2252 => x"ff2e8838",
2253 => x"74b00c87",
2254 => x"3d0d0480",
2255 => x"dfec0856",
2256 => x"75802ef0",
2257 => x"38777671",
2258 => x"0c5474b0",
2259 => x"0c873d0d",
2260 => x"04fb3d0d",
2261 => x"800b80df",
2262 => x"ec0c7a53",
2263 => x"79527851",
2264 => x"82943fb0",
2265 => x"0855b008",
2266 => x"ff2e8838",
2267 => x"74b00c87",
2268 => x"3d0d0480",
2269 => x"dfec0856",
2270 => x"75802ef0",
2271 => x"38777671",
2272 => x"0c5474b0",
2273 => x"0c873d0d",
2274 => x"04fe3d0d",
2275 => x"80dfe008",
2276 => x"51708a38",
2277 => x"80dff070",
2278 => x"80dfe00c",
2279 => x"51707512",
2280 => x"5252ff53",
2281 => x"7087fb80",
2282 => x"80268838",
2283 => x"7080dfe0",
2284 => x"0c715372",
2285 => x"b00c843d",
2286 => x"0d04fd3d",
2287 => x"0d800b80",
2288 => x"cfe40854",
2289 => x"5472812e",
2290 => x"9b387380",
2291 => x"dfe40cc2",
2292 => x"953fc0ac",
2293 => x"3f80dfb8",
2294 => x"528151c4",
2295 => x"a73fb008",
2296 => x"5185bf3f",
2297 => x"7280dfe4",
2298 => x"0cc1fb3f",
2299 => x"c0923f80",
2300 => x"dfb85281",
2301 => x"51c48d3f",
2302 => x"b0085185",
2303 => x"a53f00ff",
2304 => x"39f53d0d",
2305 => x"7e6080df",
2306 => x"e408705b",
2307 => x"585b5b75",
2308 => x"80c23877",
2309 => x"7a25a138",
2310 => x"771b7033",
2311 => x"7081ff06",
2312 => x"58585975",
2313 => x"8a2e9838",
2314 => x"7681ff06",
2315 => x"51c1963f",
2316 => x"81185879",
2317 => x"7824e138",
2318 => x"79b00c8d",
2319 => x"3d0d048d",
2320 => x"51c1823f",
2321 => x"78337081",
2322 => x"ff065257",
2323 => x"c0f73f81",
2324 => x"1858e039",
2325 => x"79557a54",
2326 => x"7d538552",
2327 => x"8d3dfc05",
2328 => x"51ffbfde",
2329 => x"3fb00856",
2330 => x"84b13f7b",
2331 => x"b0080c75",
2332 => x"b00c8d3d",
2333 => x"0d04f63d",
2334 => x"0d7d7f80",
2335 => x"dfe40870",
2336 => x"5b585a5a",
2337 => x"7580c138",
2338 => x"777925b3",
2339 => x"38c0913f",
2340 => x"b00881ff",
2341 => x"06708d32",
2342 => x"7030709f",
2343 => x"2a515157",
2344 => x"57768a2e",
2345 => x"80c43875",
2346 => x"802ebf38",
2347 => x"771a5676",
2348 => x"76347651",
2349 => x"c08f3f81",
2350 => x"18587878",
2351 => x"24cf3877",
2352 => x"5675b00c",
2353 => x"8c3d0d04",
2354 => x"78557954",
2355 => x"7c538452",
2356 => x"8c3dfc05",
2357 => x"51ffbeea",
2358 => x"3fb00856",
2359 => x"83bd3f7a",
2360 => x"b0080c75",
2361 => x"b00c8c3d",
2362 => x"0d04771a",
2363 => x"568a7634",
2364 => x"8118588d",
2365 => x"51ffbfcd",
2366 => x"3f8a51ff",
2367 => x"bfc73f77",
2368 => x"56ffbe39",
2369 => x"fb3d0d80",
2370 => x"dfe40870",
2371 => x"56547388",
2372 => x"3874b00c",
2373 => x"873d0d04",
2374 => x"77538352",
2375 => x"873dfc05",
2376 => x"51ffbe9e",
2377 => x"3fb00854",
2378 => x"82f13f75",
2379 => x"b0080c73",
2380 => x"b00c873d",
2381 => x"0d04fa3d",
2382 => x"0d80dfe4",
2383 => x"08802ea3",
2384 => x"387a5579",
2385 => x"54785386",
2386 => x"52883dfc",
2387 => x"0551ffbd",
2388 => x"f13fb008",
2389 => x"5682c43f",
2390 => x"76b0080c",
2391 => x"75b00c88",
2392 => x"3d0d0482",
2393 => x"b63f9d0b",
2394 => x"b0080cff",
2395 => x"0bb00c88",
2396 => x"3d0d04fb",
2397 => x"3d0d7779",
2398 => x"56568070",
2399 => x"54547375",
2400 => x"259f3874",
2401 => x"101010f8",
2402 => x"05527216",
2403 => x"70337074",
2404 => x"2b760781",
2405 => x"16f81656",
2406 => x"56565151",
2407 => x"747324ea",
2408 => x"3873b00c",
2409 => x"873d0d04",
2410 => x"fc3d0d76",
2411 => x"785555bc",
2412 => x"53805273",
2413 => x"51f5c63f",
2414 => x"84527451",
2415 => x"ffb53fb0",
2416 => x"08742384",
2417 => x"52841551",
2418 => x"ffa93fb0",
2419 => x"08821523",
2420 => x"84528815",
2421 => x"51ff9c3f",
2422 => x"b0088415",
2423 => x"0c84528c",
2424 => x"1551ff8f",
2425 => x"3fb00888",
2426 => x"15238452",
2427 => x"901551ff",
2428 => x"823fb008",
2429 => x"8a152384",
2430 => x"52941551",
2431 => x"fef53fb0",
2432 => x"088c1523",
2433 => x"84529815",
2434 => x"51fee83f",
2435 => x"b0088e15",
2436 => x"2388529c",
2437 => x"1551fedb",
2438 => x"3fb00890",
2439 => x"150c863d",
2440 => x"0d04e93d",
2441 => x"0d6a80df",
2442 => x"e4085757",
2443 => x"75933880",
2444 => x"c0800b84",
2445 => x"180c75ac",
2446 => x"180c75b0",
2447 => x"0c993d0d",
2448 => x"04893d70",
2449 => x"556a5455",
2450 => x"8a52993d",
2451 => x"ffbc0551",
2452 => x"ffbbef3f",
2453 => x"b0087753",
2454 => x"755256fe",
2455 => x"cb3fbc3f",
2456 => x"77b0080c",
2457 => x"75b00c99",
2458 => x"3d0d04fc",
2459 => x"3d0d8154",
2460 => x"80dfe408",
2461 => x"883873b0",
2462 => x"0c863d0d",
2463 => x"04765397",
2464 => x"b952863d",
2465 => x"fc0551ff",
2466 => x"bbb83fb0",
2467 => x"08548c3f",
2468 => x"74b0080c",
2469 => x"73b00c86",
2470 => x"3d0d0480",
2471 => x"cff408b0",
2472 => x"0c04f73d",
2473 => x"0d7b80cf",
2474 => x"f40882c8",
2475 => x"11085a54",
2476 => x"5a77802e",
2477 => x"80da3881",
2478 => x"88188419",
2479 => x"08ff0581",
2480 => x"712b5955",
2481 => x"59807424",
2482 => x"80ea3880",
2483 => x"7424b538",
2484 => x"73822b78",
2485 => x"11880556",
2486 => x"56818019",
2487 => x"08770653",
2488 => x"72802eb6",
2489 => x"38781670",
2490 => x"08535379",
2491 => x"51740853",
2492 => x"722dff14",
2493 => x"fc17fc17",
2494 => x"79812c5a",
2495 => x"57575473",
2496 => x"8025d638",
2497 => x"77085877",
2498 => x"ffad3880",
2499 => x"cff40853",
2500 => x"bc1308a5",
2501 => x"387951f9",
2502 => x"e53f7408",
2503 => x"53722dff",
2504 => x"14fc17fc",
2505 => x"1779812c",
2506 => x"5a575754",
2507 => x"738025ff",
2508 => x"a838d139",
2509 => x"8057ff93",
2510 => x"397251bc",
2511 => x"13085372",
2512 => x"2d7951f9",
2513 => x"b93fff3d",
2514 => x"0d80dfc0",
2515 => x"0bfc0570",
2516 => x"08525270",
2517 => x"ff2e9138",
2518 => x"702dfc12",
2519 => x"70085252",
2520 => x"70ff2e09",
2521 => x"8106f138",
2522 => x"833d0d04",
2523 => x"04ffbbe1",
2524 => x"3f040000",
2525 => x"00ffffff",
2526 => x"ff00ffff",
2527 => x"ffff00ff",
2528 => x"ffffff00",
2529 => x"00000040",
2530 => x"30313233",
2531 => x"34353637",
2532 => x"38396162",
2533 => x"63646566",
2534 => x"00000000",
2535 => x"2d2d0000",
2536 => x"7a776320",
2537 => x"633a0000",
2538 => x"7a776320",
2539 => x"733a0000",
2540 => x"476f7420",
2541 => x"696e7465",
2542 => x"72727570",
2543 => x"740a0000",
2544 => x"4e6f2069",
2545 => x"6e746572",
2546 => x"72757074",
2547 => x"0a000000",
2548 => x"43000000",
2549 => x"64756d6d",
2550 => x"792e6578",
2551 => x"65000000",
2552 => x"00000000",
2553 => x"00000000",
2554 => x"00000000",
2555 => x"00002fc8",
2556 => x"00002788",
2557 => x"000027f8",
2558 => x"00000000",
2559 => x"00002a60",
2560 => x"00002abc",
2561 => x"00002b18",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"00000000",
2568 => x"00000000",
2569 => x"00000000",
2570 => x"00000000",
2571 => x"000027d0",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000000",
2586 => x"00000000",
2587 => x"00000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000000",
2597 => x"00000000",
2598 => x"00000000",
2599 => x"00000000",
2600 => x"00000001",
2601 => x"330eabcd",
2602 => x"1234e66d",
2603 => x"deec0005",
2604 => x"000b0000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"ffffffff",
2794 => x"00000000",
2795 => x"00020000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00002bb0",
2799 => x"00002bb0",
2800 => x"00002bb8",
2801 => x"00002bb8",
2802 => x"00002bc0",
2803 => x"00002bc0",
2804 => x"00002bc8",
2805 => x"00002bc8",
2806 => x"00002bd0",
2807 => x"00002bd0",
2808 => x"00002bd8",
2809 => x"00002bd8",
2810 => x"00002be0",
2811 => x"00002be0",
2812 => x"00002be8",
2813 => x"00002be8",
2814 => x"00002bf0",
2815 => x"00002bf0",
2816 => x"00002bf8",
2817 => x"00002bf8",
2818 => x"00002c00",
2819 => x"00002c00",
2820 => x"00002c08",
2821 => x"00002c08",
2822 => x"00002c10",
2823 => x"00002c10",
2824 => x"00002c18",
2825 => x"00002c18",
2826 => x"00002c20",
2827 => x"00002c20",
2828 => x"00002c28",
2829 => x"00002c28",
2830 => x"00002c30",
2831 => x"00002c30",
2832 => x"00002c38",
2833 => x"00002c38",
2834 => x"00002c40",
2835 => x"00002c40",
2836 => x"00002c48",
2837 => x"00002c48",
2838 => x"00002c50",
2839 => x"00002c50",
2840 => x"00002c58",
2841 => x"00002c58",
2842 => x"00002c60",
2843 => x"00002c60",
2844 => x"00002c68",
2845 => x"00002c68",
2846 => x"00002c70",
2847 => x"00002c70",
2848 => x"00002c78",
2849 => x"00002c78",
2850 => x"00002c80",
2851 => x"00002c80",
2852 => x"00002c88",
2853 => x"00002c88",
2854 => x"00002c90",
2855 => x"00002c90",
2856 => x"00002c98",
2857 => x"00002c98",
2858 => x"00002ca0",
2859 => x"00002ca0",
2860 => x"00002ca8",
2861 => x"00002ca8",
2862 => x"00002cb0",
2863 => x"00002cb0",
2864 => x"00002cb8",
2865 => x"00002cb8",
2866 => x"00002cc0",
2867 => x"00002cc0",
2868 => x"00002cc8",
2869 => x"00002cc8",
2870 => x"00002cd0",
2871 => x"00002cd0",
2872 => x"00002cd8",
2873 => x"00002cd8",
2874 => x"00002ce0",
2875 => x"00002ce0",
2876 => x"00002ce8",
2877 => x"00002ce8",
2878 => x"00002cf0",
2879 => x"00002cf0",
2880 => x"00002cf8",
2881 => x"00002cf8",
2882 => x"00002d00",
2883 => x"00002d00",
2884 => x"00002d08",
2885 => x"00002d08",
2886 => x"00002d10",
2887 => x"00002d10",
2888 => x"00002d18",
2889 => x"00002d18",
2890 => x"00002d20",
2891 => x"00002d20",
2892 => x"00002d28",
2893 => x"00002d28",
2894 => x"00002d30",
2895 => x"00002d30",
2896 => x"00002d38",
2897 => x"00002d38",
2898 => x"00002d40",
2899 => x"00002d40",
2900 => x"00002d48",
2901 => x"00002d48",
2902 => x"00002d50",
2903 => x"00002d50",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"00002eb8",
2993 => x"00002eb8",
2994 => x"00002ec0",
2995 => x"00002ec0",
2996 => x"00002ec8",
2997 => x"00002ec8",
2998 => x"00002ed0",
2999 => x"00002ed0",
3000 => x"00002ed8",
3001 => x"00002ed8",
3002 => x"00002ee0",
3003 => x"00002ee0",
3004 => x"00002ee8",
3005 => x"00002ee8",
3006 => x"00002ef0",
3007 => x"00002ef0",
3008 => x"00002ef8",
3009 => x"00002ef8",
3010 => x"00002f00",
3011 => x"00002f00",
3012 => x"00002f08",
3013 => x"00002f08",
3014 => x"00002f10",
3015 => x"00002f10",
3016 => x"00002f18",
3017 => x"00002f18",
3018 => x"00002f20",
3019 => x"00002f20",
3020 => x"00002f28",
3021 => x"00002f28",
3022 => x"00002f30",
3023 => x"00002f30",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"00002fa0",
3051 => x"00002fa0",
3052 => x"00002fa8",
3053 => x"00002fa8",
3054 => x"000027d4",
3055 => x"ffffffff",
3056 => x"00000000",
3057 => x"ffffffff",
3058 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

