------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cdec0c",
3 => x"3a0b0b80",
4 => x"c5e80400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80cd",
162 => x"a0738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cde80c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83863f80",
257 => x"c4ec3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8d982d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8be62d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b80880c6",
294 => x"af2db80c",
295 => x"b40cb00c",
296 => x"04fe3d0d",
297 => x"0b0b80dd",
298 => x"d4085384",
299 => x"13087088",
300 => x"2a708106",
301 => x"51525270",
302 => x"802ef038",
303 => x"7181ff06",
304 => x"b00c843d",
305 => x"0d04ff3d",
306 => x"0d0b0b80",
307 => x"ddd40852",
308 => x"71087088",
309 => x"2a813270",
310 => x"81065151",
311 => x"5170f138",
312 => x"73720c83",
313 => x"3d0d0480",
314 => x"cde80880",
315 => x"2ea43880",
316 => x"cdec0882",
317 => x"2ebd3883",
318 => x"80800b0b",
319 => x"0b80ddd4",
320 => x"0c82a080",
321 => x"0b80ddd8",
322 => x"0c829080",
323 => x"0b80dddc",
324 => x"0c04f880",
325 => x"8080a40b",
326 => x"0b0b80dd",
327 => x"d40cf880",
328 => x"8082800b",
329 => x"80ddd80c",
330 => x"f8808084",
331 => x"800b80dd",
332 => x"dc0c0480",
333 => x"c0a8808c",
334 => x"0b0b0b80",
335 => x"ddd40c80",
336 => x"c0a88094",
337 => x"0b80ddd8",
338 => x"0c80cdb0",
339 => x"0b80dddc",
340 => x"0c04ff3d",
341 => x"0d80dde0",
342 => x"335170a7",
343 => x"3880cdf4",
344 => x"08700852",
345 => x"5270802e",
346 => x"94388412",
347 => x"80cdf40c",
348 => x"702d80cd",
349 => x"f4087008",
350 => x"525270ee",
351 => x"38810b80",
352 => x"dde03483",
353 => x"3d0d0404",
354 => x"803d0d0b",
355 => x"0b80ddd0",
356 => x"08802e8e",
357 => x"380b0b0b",
358 => x"0b800b80",
359 => x"2e098106",
360 => x"8538823d",
361 => x"0d040b0b",
362 => x"80ddd051",
363 => x"0b0b0bf4",
364 => x"cf3f823d",
365 => x"0d0404fe",
366 => x"3d0d8953",
367 => x"80cdb451",
368 => x"85f93f80",
369 => x"cdc45185",
370 => x"f23f810a",
371 => x"0b80ddec",
372 => x"0cff0b80",
373 => x"ddf00cff",
374 => x"13537280",
375 => x"25de3872",
376 => x"b00c843d",
377 => x"0d04bc08",
378 => x"02bc0cf9",
379 => x"3d0d800b",
380 => x"bc08fc05",
381 => x"0cbc0888",
382 => x"05088025",
383 => x"ab38bc08",
384 => x"88050830",
385 => x"bc088805",
386 => x"0c800bbc",
387 => x"08f4050c",
388 => x"bc08fc05",
389 => x"08883881",
390 => x"0bbc08f4",
391 => x"050cbc08",
392 => x"f40508bc",
393 => x"08fc050c",
394 => x"bc088c05",
395 => x"088025ab",
396 => x"38bc088c",
397 => x"050830bc",
398 => x"088c050c",
399 => x"800bbc08",
400 => x"f0050cbc",
401 => x"08fc0508",
402 => x"8838810b",
403 => x"bc08f005",
404 => x"0cbc08f0",
405 => x"0508bc08",
406 => x"fc050c80",
407 => x"53bc088c",
408 => x"050852bc",
409 => x"08880508",
410 => x"5181a73f",
411 => x"b00870bc",
412 => x"08f8050c",
413 => x"54bc08fc",
414 => x"0508802e",
415 => x"8c38bc08",
416 => x"f8050830",
417 => x"bc08f805",
418 => x"0cbc08f8",
419 => x"050870b0",
420 => x"0c54893d",
421 => x"0dbc0c04",
422 => x"bc0802bc",
423 => x"0cfb3d0d",
424 => x"800bbc08",
425 => x"fc050cbc",
426 => x"08880508",
427 => x"80259338",
428 => x"bc088805",
429 => x"0830bc08",
430 => x"88050c81",
431 => x"0bbc08fc",
432 => x"050cbc08",
433 => x"8c050880",
434 => x"258c38bc",
435 => x"088c0508",
436 => x"30bc088c",
437 => x"050c8153",
438 => x"bc088c05",
439 => x"0852bc08",
440 => x"88050851",
441 => x"ad3fb008",
442 => x"70bc08f8",
443 => x"050c54bc",
444 => x"08fc0508",
445 => x"802e8c38",
446 => x"bc08f805",
447 => x"0830bc08",
448 => x"f8050cbc",
449 => x"08f80508",
450 => x"70b00c54",
451 => x"873d0dbc",
452 => x"0c04bc08",
453 => x"02bc0cfd",
454 => x"3d0d810b",
455 => x"bc08fc05",
456 => x"0c800bbc",
457 => x"08f8050c",
458 => x"bc088c05",
459 => x"08bc0888",
460 => x"050827ac",
461 => x"38bc08fc",
462 => x"0508802e",
463 => x"a338800b",
464 => x"bc088c05",
465 => x"08249938",
466 => x"bc088c05",
467 => x"0810bc08",
468 => x"8c050cbc",
469 => x"08fc0508",
470 => x"10bc08fc",
471 => x"050cc939",
472 => x"bc08fc05",
473 => x"08802e80",
474 => x"c938bc08",
475 => x"8c0508bc",
476 => x"08880508",
477 => x"26a138bc",
478 => x"08880508",
479 => x"bc088c05",
480 => x"0831bc08",
481 => x"88050cbc",
482 => x"08f80508",
483 => x"bc08fc05",
484 => x"0807bc08",
485 => x"f8050cbc",
486 => x"08fc0508",
487 => x"812abc08",
488 => x"fc050cbc",
489 => x"088c0508",
490 => x"812abc08",
491 => x"8c050cff",
492 => x"af39bc08",
493 => x"90050880",
494 => x"2e8f38bc",
495 => x"08880508",
496 => x"70bc08f4",
497 => x"050c518d",
498 => x"39bc08f8",
499 => x"050870bc",
500 => x"08f4050c",
501 => x"51bc08f4",
502 => x"0508b00c",
503 => x"853d0dbc",
504 => x"0c04fc3d",
505 => x"0d767079",
506 => x"7b555555",
507 => x"558f7227",
508 => x"8c387275",
509 => x"07830651",
510 => x"70802ea7",
511 => x"38ff1252",
512 => x"71ff2e98",
513 => x"38727081",
514 => x"05543374",
515 => x"70810556",
516 => x"34ff1252",
517 => x"71ff2e09",
518 => x"8106ea38",
519 => x"74b00c86",
520 => x"3d0d0474",
521 => x"51727084",
522 => x"05540871",
523 => x"70840553",
524 => x"0c727084",
525 => x"05540871",
526 => x"70840553",
527 => x"0c727084",
528 => x"05540871",
529 => x"70840553",
530 => x"0c727084",
531 => x"05540871",
532 => x"70840553",
533 => x"0cf01252",
534 => x"718f26c9",
535 => x"38837227",
536 => x"95387270",
537 => x"84055408",
538 => x"71708405",
539 => x"530cfc12",
540 => x"52718326",
541 => x"ed387054",
542 => x"ff8339f7",
543 => x"3d0d7c70",
544 => x"525380c8",
545 => x"3f7254b0",
546 => x"085580cd",
547 => x"d4568157",
548 => x"b0088105",
549 => x"5a8b3de4",
550 => x"11595382",
551 => x"59f41352",
552 => x"7b881108",
553 => x"52538183",
554 => x"3fb00830",
555 => x"70b00807",
556 => x"9f2c8a07",
557 => x"b00c538b",
558 => x"3d0d04ff",
559 => x"3d0d7352",
560 => x"80cdf808",
561 => x"51ffb43f",
562 => x"833d0d04",
563 => x"fd3d0d75",
564 => x"70718306",
565 => x"53555270",
566 => x"b8387170",
567 => x"087009f7",
568 => x"fbfdff12",
569 => x"0670f884",
570 => x"82818006",
571 => x"51515253",
572 => x"709d3884",
573 => x"13700870",
574 => x"09f7fbfd",
575 => x"ff120670",
576 => x"f8848281",
577 => x"80065151",
578 => x"52537080",
579 => x"2ee53872",
580 => x"52713351",
581 => x"70802e8a",
582 => x"38811270",
583 => x"33525270",
584 => x"f8387174",
585 => x"31b00c85",
586 => x"3d0d04f2",
587 => x"3d0d6062",
588 => x"88110870",
589 => x"57575f5a",
590 => x"74802e81",
591 => x"8f388c1a",
592 => x"2270832a",
593 => x"81327081",
594 => x"06515558",
595 => x"73863890",
596 => x"1a089138",
597 => x"795190a1",
598 => x"3fff54b0",
599 => x"0880ed38",
600 => x"8c1a2258",
601 => x"7d085780",
602 => x"7883ffff",
603 => x"0670812a",
604 => x"70810651",
605 => x"56575573",
606 => x"752e80d7",
607 => x"38749038",
608 => x"76088418",
609 => x"08881959",
610 => x"56597480",
611 => x"2ef23874",
612 => x"54888075",
613 => x"27843888",
614 => x"80547353",
615 => x"78529c1a",
616 => x"0851a41a",
617 => x"0854732d",
618 => x"800bb008",
619 => x"2582e638",
620 => x"b0081975",
621 => x"b008317f",
622 => x"880508b0",
623 => x"08317061",
624 => x"88050c56",
625 => x"565973ff",
626 => x"b4388054",
627 => x"73b00c90",
628 => x"3d0d0475",
629 => x"81327081",
630 => x"06764151",
631 => x"5473802e",
632 => x"81c13874",
633 => x"90387608",
634 => x"84180888",
635 => x"19595659",
636 => x"74802ef2",
637 => x"38881a08",
638 => x"7883ffff",
639 => x"0670892a",
640 => x"70810651",
641 => x"56595673",
642 => x"802e82fa",
643 => x"38757527",
644 => x"8d387787",
645 => x"2a708106",
646 => x"51547382",
647 => x"b5387476",
648 => x"27833874",
649 => x"56755378",
650 => x"52790851",
651 => x"85823f88",
652 => x"1a087631",
653 => x"881b0c79",
654 => x"08167a0c",
655 => x"74567519",
656 => x"7577317f",
657 => x"88050878",
658 => x"31706188",
659 => x"050c5656",
660 => x"5973802e",
661 => x"fef4388c",
662 => x"1a2258ff",
663 => x"86397778",
664 => x"5479537b",
665 => x"525684c8",
666 => x"3f881a08",
667 => x"7831881b",
668 => x"0c790818",
669 => x"7a0c7c76",
670 => x"315d7c8e",
671 => x"3879518f",
672 => x"db3fb008",
673 => x"818f38b0",
674 => x"085f7519",
675 => x"7577317f",
676 => x"88050878",
677 => x"31706188",
678 => x"050c5656",
679 => x"5973802e",
680 => x"fea83874",
681 => x"81833876",
682 => x"08841808",
683 => x"88195956",
684 => x"5974802e",
685 => x"f2387453",
686 => x"8a527851",
687 => x"82d33fb0",
688 => x"08793181",
689 => x"055db008",
690 => x"84388115",
691 => x"5d815f7c",
692 => x"58747d27",
693 => x"83387458",
694 => x"941a0888",
695 => x"1b081157",
696 => x"5c807a08",
697 => x"5c54901a",
698 => x"087b2783",
699 => x"38815475",
700 => x"78258438",
701 => x"73ba387b",
702 => x"7824fee2",
703 => x"387b5378",
704 => x"529c1a08",
705 => x"51a41a08",
706 => x"54732db0",
707 => x"0856b008",
708 => x"8024fee2",
709 => x"388c1a22",
710 => x"80c00754",
711 => x"738c1b23",
712 => x"ff5473b0",
713 => x"0c903d0d",
714 => x"047effa3",
715 => x"38ff8739",
716 => x"75537852",
717 => x"7a5182f8",
718 => x"3f790816",
719 => x"7a0c7951",
720 => x"8e9a3fb0",
721 => x"08cf387c",
722 => x"76315d7c",
723 => x"febc38fe",
724 => x"ac39901a",
725 => x"087a0871",
726 => x"31761170",
727 => x"565a5752",
728 => x"80cdf808",
729 => x"51848c3f",
730 => x"b008802e",
731 => x"ffa738b0",
732 => x"08901b0c",
733 => x"b008167a",
734 => x"0c77941b",
735 => x"0c74881b",
736 => x"0c7456fd",
737 => x"99397908",
738 => x"58901a08",
739 => x"78278338",
740 => x"81547575",
741 => x"27843873",
742 => x"b338941a",
743 => x"08567575",
744 => x"2680d338",
745 => x"75537852",
746 => x"9c1a0851",
747 => x"a41a0854",
748 => x"732db008",
749 => x"56b00880",
750 => x"24fd8338",
751 => x"8c1a2280",
752 => x"c0075473",
753 => x"8c1b23ff",
754 => x"54fed739",
755 => x"75537852",
756 => x"775181dc",
757 => x"3f790816",
758 => x"7a0c7951",
759 => x"8cfe3fb0",
760 => x"08802efc",
761 => x"d9388c1a",
762 => x"2280c007",
763 => x"54738c1b",
764 => x"23ff54fe",
765 => x"ad397475",
766 => x"54795378",
767 => x"525681b0",
768 => x"3f881a08",
769 => x"7531881b",
770 => x"0c790815",
771 => x"7a0cfcae",
772 => x"39fa3d0d",
773 => x"7a790288",
774 => x"05a70533",
775 => x"56525383",
776 => x"73278a38",
777 => x"70830652",
778 => x"71802ea8",
779 => x"38ff1353",
780 => x"72ff2e97",
781 => x"38703352",
782 => x"73722e91",
783 => x"388111ff",
784 => x"14545172",
785 => x"ff2e0981",
786 => x"06eb3880",
787 => x"5170b00c",
788 => x"883d0d04",
789 => x"70725755",
790 => x"83517582",
791 => x"802914ff",
792 => x"12525670",
793 => x"8025f338",
794 => x"837327bf",
795 => x"38740876",
796 => x"327009f7",
797 => x"fbfdff12",
798 => x"0670f884",
799 => x"82818006",
800 => x"51515170",
801 => x"802e9938",
802 => x"74518052",
803 => x"70335773",
804 => x"772effb9",
805 => x"38811181",
806 => x"13535183",
807 => x"7227ed38",
808 => x"fc138416",
809 => x"56537283",
810 => x"26c33874",
811 => x"51fefe39",
812 => x"fa3d0d78",
813 => x"7a7c7272",
814 => x"72575757",
815 => x"59565674",
816 => x"7627b238",
817 => x"76155175",
818 => x"7127aa38",
819 => x"707717ff",
820 => x"14545553",
821 => x"71ff2e96",
822 => x"38ff14ff",
823 => x"14545472",
824 => x"337434ff",
825 => x"125271ff",
826 => x"2e098106",
827 => x"ec3875b0",
828 => x"0c883d0d",
829 => x"04768f26",
830 => x"9738ff12",
831 => x"5271ff2e",
832 => x"ed387270",
833 => x"81055433",
834 => x"74708105",
835 => x"5634eb39",
836 => x"74760783",
837 => x"065170e2",
838 => x"38757554",
839 => x"51727084",
840 => x"05540871",
841 => x"70840553",
842 => x"0c727084",
843 => x"05540871",
844 => x"70840553",
845 => x"0c727084",
846 => x"05540871",
847 => x"70840553",
848 => x"0c727084",
849 => x"05540871",
850 => x"70840553",
851 => x"0cf01252",
852 => x"718f26c9",
853 => x"38837227",
854 => x"95387270",
855 => x"84055408",
856 => x"71708405",
857 => x"530cfc12",
858 => x"52718326",
859 => x"ed387054",
860 => x"ff8839ef",
861 => x"3d0d6365",
862 => x"67405d42",
863 => x"7b802e84",
864 => x"fa386151",
865 => x"a5b43ff8",
866 => x"1c708412",
867 => x"0870fc06",
868 => x"70628b05",
869 => x"70f80641",
870 => x"59455b5c",
871 => x"41579674",
872 => x"2782c338",
873 => x"807b247e",
874 => x"7c260759",
875 => x"80547874",
876 => x"2e098106",
877 => x"82a93877",
878 => x"7b2581fc",
879 => x"38771780",
880 => x"d5b40b88",
881 => x"05085e56",
882 => x"7c762e84",
883 => x"bd388416",
884 => x"0870fe06",
885 => x"17841108",
886 => x"81065155",
887 => x"5573828b",
888 => x"3874fc06",
889 => x"597c762e",
890 => x"84dd3877",
891 => x"195f7e7b",
892 => x"2581fd38",
893 => x"79810654",
894 => x"7382bf38",
895 => x"76770831",
896 => x"841108fc",
897 => x"06565a75",
898 => x"802e9138",
899 => x"7c762e84",
900 => x"ea387419",
901 => x"1859787b",
902 => x"25848938",
903 => x"79802e82",
904 => x"99387715",
905 => x"567a7624",
906 => x"8290388c",
907 => x"1a08881b",
908 => x"08718c12",
909 => x"0c88120c",
910 => x"55797659",
911 => x"57881761",
912 => x"fc055759",
913 => x"75a42685",
914 => x"ef387b79",
915 => x"55559376",
916 => x"2780c938",
917 => x"7b708405",
918 => x"5d087c56",
919 => x"790c7470",
920 => x"84055608",
921 => x"8c180c90",
922 => x"17549b76",
923 => x"27ae3874",
924 => x"70840556",
925 => x"08740c74",
926 => x"70840556",
927 => x"0894180c",
928 => x"981754a3",
929 => x"76279538",
930 => x"74708405",
931 => x"5608740c",
932 => x"74708405",
933 => x"56089c18",
934 => x"0ca01754",
935 => x"74708405",
936 => x"56087470",
937 => x"8405560c",
938 => x"74708405",
939 => x"56087470",
940 => x"8405560c",
941 => x"7408740c",
942 => x"777b3156",
943 => x"758f2680",
944 => x"c9388417",
945 => x"08810678",
946 => x"0784180c",
947 => x"77178411",
948 => x"08810784",
949 => x"120c5461",
950 => x"51a2e03f",
951 => x"88175473",
952 => x"b00c933d",
953 => x"0d04905b",
954 => x"fdba3978",
955 => x"56fe8539",
956 => x"8c160888",
957 => x"1708718c",
958 => x"120c8812",
959 => x"0c557e70",
960 => x"7c315758",
961 => x"8f7627ff",
962 => x"b9387a17",
963 => x"84180881",
964 => x"067c0784",
965 => x"190c7681",
966 => x"0784120c",
967 => x"76118411",
968 => x"08810784",
969 => x"120c5588",
970 => x"05526151",
971 => x"8cf63f61",
972 => x"51a2883f",
973 => x"881754ff",
974 => x"a6397d52",
975 => x"615194f5",
976 => x"3fb00859",
977 => x"b008802e",
978 => x"81a338b0",
979 => x"08f80560",
980 => x"840508fe",
981 => x"06610555",
982 => x"5776742e",
983 => x"83e638fc",
984 => x"185675a4",
985 => x"2681aa38",
986 => x"7bb00855",
987 => x"55937627",
988 => x"80d83874",
989 => x"70840556",
990 => x"08b00870",
991 => x"8405b00c",
992 => x"0cb00875",
993 => x"70840557",
994 => x"08717084",
995 => x"05530c54",
996 => x"9b7627b6",
997 => x"38747084",
998 => x"05560874",
999 => x"70840556",
1000 => x"0c747084",
1001 => x"05560874",
1002 => x"70840556",
1003 => x"0ca37627",
1004 => x"99387470",
1005 => x"84055608",
1006 => x"74708405",
1007 => x"560c7470",
1008 => x"84055608",
1009 => x"74708405",
1010 => x"560c7470",
1011 => x"84055608",
1012 => x"74708405",
1013 => x"560c7470",
1014 => x"84055608",
1015 => x"74708405",
1016 => x"560c7408",
1017 => x"740c7b52",
1018 => x"61518bb8",
1019 => x"3f6151a0",
1020 => x"ca3f7854",
1021 => x"73b00c93",
1022 => x"3d0d047d",
1023 => x"52615193",
1024 => x"b43fb008",
1025 => x"b00c933d",
1026 => x"0d048416",
1027 => x"0855fbd1",
1028 => x"3975537b",
1029 => x"52b00851",
1030 => x"efc83f7b",
1031 => x"5261518b",
1032 => x"833fca39",
1033 => x"8c160888",
1034 => x"1708718c",
1035 => x"120c8812",
1036 => x"0c558c1a",
1037 => x"08881b08",
1038 => x"718c120c",
1039 => x"88120c55",
1040 => x"79795957",
1041 => x"fbf73977",
1042 => x"19901c55",
1043 => x"55737524",
1044 => x"fba2387a",
1045 => x"177080d5",
1046 => x"b40b8805",
1047 => x"0c757c31",
1048 => x"81078412",
1049 => x"0c5d8417",
1050 => x"0881067b",
1051 => x"0784180c",
1052 => x"61519fc7",
1053 => x"3f881754",
1054 => x"fce53974",
1055 => x"1918901c",
1056 => x"555d737d",
1057 => x"24fb9538",
1058 => x"8c1a0888",
1059 => x"1b08718c",
1060 => x"120c8812",
1061 => x"0c55881a",
1062 => x"61fc0557",
1063 => x"5975a426",
1064 => x"81ae387b",
1065 => x"79555593",
1066 => x"762780c9",
1067 => x"387b7084",
1068 => x"055d087c",
1069 => x"56790c74",
1070 => x"70840556",
1071 => x"088c1b0c",
1072 => x"901a549b",
1073 => x"7627ae38",
1074 => x"74708405",
1075 => x"5608740c",
1076 => x"74708405",
1077 => x"5608941b",
1078 => x"0c981a54",
1079 => x"a3762795",
1080 => x"38747084",
1081 => x"05560874",
1082 => x"0c747084",
1083 => x"0556089c",
1084 => x"1b0ca01a",
1085 => x"54747084",
1086 => x"05560874",
1087 => x"70840556",
1088 => x"0c747084",
1089 => x"05560874",
1090 => x"70840556",
1091 => x"0c740874",
1092 => x"0c7a1a70",
1093 => x"80d5b40b",
1094 => x"88050c7d",
1095 => x"7c318107",
1096 => x"84120c54",
1097 => x"841a0881",
1098 => x"067b0784",
1099 => x"1b0c6151",
1100 => x"9e893f78",
1101 => x"54fdbd39",
1102 => x"75537b52",
1103 => x"7851eda2",
1104 => x"3ffaf539",
1105 => x"841708fc",
1106 => x"06186058",
1107 => x"58fae939",
1108 => x"75537b52",
1109 => x"7851ed8a",
1110 => x"3f7a1a70",
1111 => x"80d5b40b",
1112 => x"88050c7d",
1113 => x"7c318107",
1114 => x"84120c54",
1115 => x"841a0881",
1116 => x"067b0784",
1117 => x"1b0cffb6",
1118 => x"39fa3d0d",
1119 => x"7880cdf8",
1120 => x"085455b8",
1121 => x"1308802e",
1122 => x"81b5388c",
1123 => x"15227083",
1124 => x"ffff0670",
1125 => x"832a8132",
1126 => x"70810651",
1127 => x"55555672",
1128 => x"802e80dc",
1129 => x"3873842a",
1130 => x"81328106",
1131 => x"57ff5376",
1132 => x"80f63873",
1133 => x"822a7081",
1134 => x"06515372",
1135 => x"802eb938",
1136 => x"b0150854",
1137 => x"73802e9c",
1138 => x"3880c015",
1139 => x"5373732e",
1140 => x"8f387352",
1141 => x"80cdf808",
1142 => x"5187c93f",
1143 => x"8c152256",
1144 => x"76b0160c",
1145 => x"75db0653",
1146 => x"728c1623",
1147 => x"800b8416",
1148 => x"0c901508",
1149 => x"750c7256",
1150 => x"75880753",
1151 => x"728c1623",
1152 => x"90150880",
1153 => x"2e80c038",
1154 => x"8c152270",
1155 => x"81065553",
1156 => x"739d3872",
1157 => x"812a7081",
1158 => x"06515372",
1159 => x"85389415",
1160 => x"08547388",
1161 => x"160c8053",
1162 => x"72b00c88",
1163 => x"3d0d0480",
1164 => x"0b88160c",
1165 => x"94150830",
1166 => x"98160c80",
1167 => x"53ea3972",
1168 => x"5182fb3f",
1169 => x"fec53974",
1170 => x"518ce83f",
1171 => x"8c152270",
1172 => x"81065553",
1173 => x"73802eff",
1174 => x"ba38d439",
1175 => x"f83d0d7a",
1176 => x"5877802e",
1177 => x"81993880",
1178 => x"cdf80854",
1179 => x"b8140880",
1180 => x"2e80ed38",
1181 => x"8c182270",
1182 => x"902b7090",
1183 => x"2c70832a",
1184 => x"81328106",
1185 => x"5c515754",
1186 => x"7880cd38",
1187 => x"90180857",
1188 => x"76802e80",
1189 => x"c3387708",
1190 => x"77317779",
1191 => x"0c768306",
1192 => x"7a585555",
1193 => x"73853894",
1194 => x"18085675",
1195 => x"88190c80",
1196 => x"7525a538",
1197 => x"74537652",
1198 => x"9c180851",
1199 => x"a4180854",
1200 => x"732d800b",
1201 => x"b0082580",
1202 => x"c938b008",
1203 => x"1775b008",
1204 => x"31565774",
1205 => x"8024dd38",
1206 => x"800bb00c",
1207 => x"8a3d0d04",
1208 => x"735181da",
1209 => x"3f8c1822",
1210 => x"70902b70",
1211 => x"902c7083",
1212 => x"2a813281",
1213 => x"065c5157",
1214 => x"5478dd38",
1215 => x"ff8e39a4",
1216 => x"dc5280cd",
1217 => x"f8085189",
1218 => x"f13fb008",
1219 => x"b00c8a3d",
1220 => x"0d048c18",
1221 => x"2280c007",
1222 => x"54738c19",
1223 => x"23ff0bb0",
1224 => x"0c8a3d0d",
1225 => x"04803d0d",
1226 => x"72518071",
1227 => x"0c800b84",
1228 => x"120c800b",
1229 => x"88120c02",
1230 => x"8e05228c",
1231 => x"12230292",
1232 => x"05228e12",
1233 => x"23800b90",
1234 => x"120c800b",
1235 => x"94120c80",
1236 => x"0b98120c",
1237 => x"709c120c",
1238 => x"80c0f00b",
1239 => x"a0120c80",
1240 => x"c1bc0ba4",
1241 => x"120c80c2",
1242 => x"b80ba812",
1243 => x"0c80c389",
1244 => x"0bac120c",
1245 => x"823d0d04",
1246 => x"fa3d0d79",
1247 => x"7080dc29",
1248 => x"8c11547a",
1249 => x"5356578c",
1250 => x"ac3fb008",
1251 => x"b0085556",
1252 => x"b008802e",
1253 => x"a238b008",
1254 => x"8c055480",
1255 => x"0bb0080c",
1256 => x"76b00884",
1257 => x"050c73b0",
1258 => x"0888050c",
1259 => x"74538052",
1260 => x"735197f7",
1261 => x"3f755473",
1262 => x"b00c883d",
1263 => x"0d04fc3d",
1264 => x"0d76a9d1",
1265 => x"0bbc120c",
1266 => x"55810bb8",
1267 => x"160c800b",
1268 => x"84dc160c",
1269 => x"830b84e0",
1270 => x"160c84e8",
1271 => x"1584e416",
1272 => x"0c745480",
1273 => x"53845284",
1274 => x"150851fe",
1275 => x"b83f7454",
1276 => x"81538952",
1277 => x"88150851",
1278 => x"feab3f74",
1279 => x"5482538a",
1280 => x"528c1508",
1281 => x"51fe9e3f",
1282 => x"863d0d04",
1283 => x"f93d0d79",
1284 => x"80cdf808",
1285 => x"5457b813",
1286 => x"08802e80",
1287 => x"c83884dc",
1288 => x"13568816",
1289 => x"08841708",
1290 => x"ff055555",
1291 => x"8074249f",
1292 => x"388c1522",
1293 => x"70902b70",
1294 => x"902c5154",
1295 => x"5872802e",
1296 => x"80ca3880",
1297 => x"dc15ff15",
1298 => x"55557380",
1299 => x"25e33875",
1300 => x"08537280",
1301 => x"2e9f3872",
1302 => x"56881608",
1303 => x"841708ff",
1304 => x"055555c8",
1305 => x"397251fe",
1306 => x"d53f80cd",
1307 => x"f80884dc",
1308 => x"0556ffae",
1309 => x"39845276",
1310 => x"51fdfd3f",
1311 => x"b008760c",
1312 => x"b008802e",
1313 => x"80c038b0",
1314 => x"0856ce39",
1315 => x"810b8c16",
1316 => x"2372750c",
1317 => x"7288160c",
1318 => x"7284160c",
1319 => x"7290160c",
1320 => x"7294160c",
1321 => x"7298160c",
1322 => x"ff0b8e16",
1323 => x"2372b016",
1324 => x"0c72b416",
1325 => x"0c7280c4",
1326 => x"160c7280",
1327 => x"c8160c74",
1328 => x"b00c893d",
1329 => x"0d048c77",
1330 => x"0c800bb0",
1331 => x"0c893d0d",
1332 => x"04ff3d0d",
1333 => x"a4dc5273",
1334 => x"51869f3f",
1335 => x"833d0d04",
1336 => x"803d0d80",
1337 => x"cdf80851",
1338 => x"e83f823d",
1339 => x"0d04fb3d",
1340 => x"0d777052",
1341 => x"5696c33f",
1342 => x"80d5b40b",
1343 => x"88050884",
1344 => x"1108fc06",
1345 => x"707b319f",
1346 => x"ef05e080",
1347 => x"06e08005",
1348 => x"565653a0",
1349 => x"80742494",
1350 => x"38805275",
1351 => x"51969d3f",
1352 => x"80d5bc08",
1353 => x"155372b0",
1354 => x"082e8f38",
1355 => x"7551968b",
1356 => x"3f805372",
1357 => x"b00c873d",
1358 => x"0d047330",
1359 => x"52755195",
1360 => x"fb3fb008",
1361 => x"ff2ea838",
1362 => x"80d5b40b",
1363 => x"88050875",
1364 => x"75318107",
1365 => x"84120c53",
1366 => x"80d4f808",
1367 => x"743180d4",
1368 => x"f80c7551",
1369 => x"95d53f81",
1370 => x"0bb00c87",
1371 => x"3d0d0480",
1372 => x"52755195",
1373 => x"c73f80d5",
1374 => x"b40b8805",
1375 => x"08b00871",
1376 => x"3156538f",
1377 => x"7525ffa4",
1378 => x"38b00880",
1379 => x"d5a80831",
1380 => x"80d4f80c",
1381 => x"74810784",
1382 => x"140c7551",
1383 => x"959d3f80",
1384 => x"53ff9039",
1385 => x"f63d0d7c",
1386 => x"7e545b72",
1387 => x"802e8283",
1388 => x"387a5195",
1389 => x"853ff813",
1390 => x"84110870",
1391 => x"fe067013",
1392 => x"841108fc",
1393 => x"065d5859",
1394 => x"545880d5",
1395 => x"bc08752e",
1396 => x"82de3878",
1397 => x"84160c80",
1398 => x"73810654",
1399 => x"5a727a2e",
1400 => x"81d53878",
1401 => x"15841108",
1402 => x"81065153",
1403 => x"72a03878",
1404 => x"17577981",
1405 => x"e6388815",
1406 => x"08537280",
1407 => x"d5bc2e82",
1408 => x"f9388c15",
1409 => x"08708c15",
1410 => x"0c738812",
1411 => x"0c567681",
1412 => x"0784190c",
1413 => x"76187771",
1414 => x"0c537981",
1415 => x"913883ff",
1416 => x"772781c8",
1417 => x"3876892a",
1418 => x"77832a56",
1419 => x"5372802e",
1420 => x"bf387686",
1421 => x"2ab80555",
1422 => x"847327b4",
1423 => x"3880db13",
1424 => x"55947327",
1425 => x"ab38768c",
1426 => x"2a80ee05",
1427 => x"5580d473",
1428 => x"279e3876",
1429 => x"8f2a80f7",
1430 => x"055582d4",
1431 => x"73279138",
1432 => x"76922a80",
1433 => x"fc05558a",
1434 => x"d4732784",
1435 => x"3880fe55",
1436 => x"74101010",
1437 => x"80d5b405",
1438 => x"88110855",
1439 => x"5673762e",
1440 => x"82b33884",
1441 => x"1408fc06",
1442 => x"53767327",
1443 => x"8d388814",
1444 => x"08547376",
1445 => x"2e098106",
1446 => x"ea388c14",
1447 => x"08708c1a",
1448 => x"0c74881a",
1449 => x"0c788812",
1450 => x"0c56778c",
1451 => x"150c7a51",
1452 => x"93893f8c",
1453 => x"3d0d0477",
1454 => x"08787131",
1455 => x"59770588",
1456 => x"19085457",
1457 => x"7280d5bc",
1458 => x"2e80e038",
1459 => x"8c180870",
1460 => x"8c150c73",
1461 => x"88120c56",
1462 => x"fe893988",
1463 => x"15088c16",
1464 => x"08708c13",
1465 => x"0c578817",
1466 => x"0cfea339",
1467 => x"76832a70",
1468 => x"54558075",
1469 => x"24819838",
1470 => x"72822c81",
1471 => x"712b80d5",
1472 => x"b8080780",
1473 => x"d5b40b84",
1474 => x"050c5374",
1475 => x"10101080",
1476 => x"d5b40588",
1477 => x"11085556",
1478 => x"758c190c",
1479 => x"7388190c",
1480 => x"7788170c",
1481 => x"778c150c",
1482 => x"ff843981",
1483 => x"5afdb439",
1484 => x"78177381",
1485 => x"06545772",
1486 => x"98387708",
1487 => x"78713159",
1488 => x"77058c19",
1489 => x"08881a08",
1490 => x"718c120c",
1491 => x"88120c57",
1492 => x"57768107",
1493 => x"84190c77",
1494 => x"80d5b40b",
1495 => x"88050c80",
1496 => x"d5b00877",
1497 => x"26fec738",
1498 => x"80d5ac08",
1499 => x"527a51fa",
1500 => x"fd3f7a51",
1501 => x"91c53ffe",
1502 => x"ba398178",
1503 => x"8c150c78",
1504 => x"88150c73",
1505 => x"8c1a0c73",
1506 => x"881a0c5a",
1507 => x"fd803983",
1508 => x"1570822c",
1509 => x"81712b80",
1510 => x"d5b80807",
1511 => x"80d5b40b",
1512 => x"84050c51",
1513 => x"53741010",
1514 => x"1080d5b4",
1515 => x"05881108",
1516 => x"5556fee4",
1517 => x"39745380",
1518 => x"7524a738",
1519 => x"72822c81",
1520 => x"712b80d5",
1521 => x"b8080780",
1522 => x"d5b40b84",
1523 => x"050c5375",
1524 => x"8c190c73",
1525 => x"88190c77",
1526 => x"88170c77",
1527 => x"8c150cfd",
1528 => x"cd398315",
1529 => x"70822c81",
1530 => x"712b80d5",
1531 => x"b8080780",
1532 => x"d5b40b84",
1533 => x"050c5153",
1534 => x"d639f93d",
1535 => x"0d797b58",
1536 => x"53800b80",
1537 => x"cdf80853",
1538 => x"5672722e",
1539 => x"80c03884",
1540 => x"dc135574",
1541 => x"762eb738",
1542 => x"88150884",
1543 => x"1608ff05",
1544 => x"54548073",
1545 => x"249d388c",
1546 => x"14227090",
1547 => x"2b70902c",
1548 => x"51535871",
1549 => x"80d83880",
1550 => x"dc14ff14",
1551 => x"54547280",
1552 => x"25e53874",
1553 => x"085574d0",
1554 => x"3880cdf8",
1555 => x"085284dc",
1556 => x"12557480",
1557 => x"2eb13888",
1558 => x"15088416",
1559 => x"08ff0554",
1560 => x"54807324",
1561 => x"9c388c14",
1562 => x"2270902b",
1563 => x"70902c51",
1564 => x"535871ad",
1565 => x"3880dc14",
1566 => x"ff145454",
1567 => x"728025e6",
1568 => x"38740855",
1569 => x"74d13875",
1570 => x"b00c893d",
1571 => x"0d047351",
1572 => x"762d75b0",
1573 => x"080780dc",
1574 => x"15ff1555",
1575 => x"5556ff9e",
1576 => x"39735176",
1577 => x"2d75b008",
1578 => x"0780dc15",
1579 => x"ff155555",
1580 => x"56ca39ea",
1581 => x"3d0d688c",
1582 => x"11227081",
1583 => x"2a810657",
1584 => x"58567480",
1585 => x"e4388e16",
1586 => x"2270902b",
1587 => x"70902c51",
1588 => x"55588074",
1589 => x"24b13898",
1590 => x"3dc40553",
1591 => x"735280cd",
1592 => x"f8085192",
1593 => x"ac3f800b",
1594 => x"b0082497",
1595 => x"387983e0",
1596 => x"80065473",
1597 => x"80c0802e",
1598 => x"818f3873",
1599 => x"8280802e",
1600 => x"8191388c",
1601 => x"16225776",
1602 => x"90800754",
1603 => x"738c1723",
1604 => x"88805280",
1605 => x"cdf80851",
1606 => x"819b3fb0",
1607 => x"089d388c",
1608 => x"16228207",
1609 => x"54738c17",
1610 => x"2380c316",
1611 => x"70770c90",
1612 => x"170c810b",
1613 => x"94170c98",
1614 => x"3d0d0480",
1615 => x"cdf808a9",
1616 => x"d10bbc12",
1617 => x"0c548c16",
1618 => x"22818007",
1619 => x"54738c17",
1620 => x"23b00876",
1621 => x"0cb00890",
1622 => x"170c8880",
1623 => x"0b94170c",
1624 => x"74802ed3",
1625 => x"388e1622",
1626 => x"70902b70",
1627 => x"902c5355",
1628 => x"5898a43f",
1629 => x"b008802e",
1630 => x"ffbd388c",
1631 => x"16228107",
1632 => x"54738c17",
1633 => x"23983d0d",
1634 => x"04810b8c",
1635 => x"17225855",
1636 => x"fef539a8",
1637 => x"160880c2",
1638 => x"b82e0981",
1639 => x"06fee438",
1640 => x"8c162288",
1641 => x"80075473",
1642 => x"8c172388",
1643 => x"800b80cc",
1644 => x"170cfedc",
1645 => x"39f33d0d",
1646 => x"7f618b11",
1647 => x"70f8065c",
1648 => x"55555e72",
1649 => x"96268338",
1650 => x"90598079",
1651 => x"24747a26",
1652 => x"07538054",
1653 => x"72742e09",
1654 => x"810680cb",
1655 => x"387d518c",
1656 => x"d93f7883",
1657 => x"f72680c6",
1658 => x"3878832a",
1659 => x"70101010",
1660 => x"80d5b405",
1661 => x"8c110859",
1662 => x"595a7678",
1663 => x"2e83b038",
1664 => x"841708fc",
1665 => x"06568c17",
1666 => x"08881808",
1667 => x"718c120c",
1668 => x"88120c58",
1669 => x"75178411",
1670 => x"08810784",
1671 => x"120c537d",
1672 => x"518c983f",
1673 => x"88175473",
1674 => x"b00c8f3d",
1675 => x"0d047889",
1676 => x"2a79832a",
1677 => x"5b537280",
1678 => x"2ebf3878",
1679 => x"862ab805",
1680 => x"5a847327",
1681 => x"b43880db",
1682 => x"135a9473",
1683 => x"27ab3878",
1684 => x"8c2a80ee",
1685 => x"055a80d4",
1686 => x"73279e38",
1687 => x"788f2a80",
1688 => x"f7055a82",
1689 => x"d4732791",
1690 => x"3878922a",
1691 => x"80fc055a",
1692 => x"8ad47327",
1693 => x"843880fe",
1694 => x"5a791010",
1695 => x"1080d5b4",
1696 => x"058c1108",
1697 => x"58557675",
1698 => x"2ea33884",
1699 => x"1708fc06",
1700 => x"707a3155",
1701 => x"56738f24",
1702 => x"88d53873",
1703 => x"8025fee6",
1704 => x"388c1708",
1705 => x"5776752e",
1706 => x"098106df",
1707 => x"38811a5a",
1708 => x"80d5c408",
1709 => x"577680d5",
1710 => x"bc2e82c0",
1711 => x"38841708",
1712 => x"fc06707a",
1713 => x"31555673",
1714 => x"8f2481f9",
1715 => x"3880d5bc",
1716 => x"0b80d5c8",
1717 => x"0c80d5bc",
1718 => x"0b80d5c4",
1719 => x"0c738025",
1720 => x"feb23883",
1721 => x"ff762783",
1722 => x"df387589",
1723 => x"2a76832a",
1724 => x"55537280",
1725 => x"2ebf3875",
1726 => x"862ab805",
1727 => x"54847327",
1728 => x"b43880db",
1729 => x"13549473",
1730 => x"27ab3875",
1731 => x"8c2a80ee",
1732 => x"055480d4",
1733 => x"73279e38",
1734 => x"758f2a80",
1735 => x"f7055482",
1736 => x"d4732791",
1737 => x"3875922a",
1738 => x"80fc0554",
1739 => x"8ad47327",
1740 => x"843880fe",
1741 => x"54731010",
1742 => x"1080d5b4",
1743 => x"05881108",
1744 => x"56587478",
1745 => x"2e86cf38",
1746 => x"841508fc",
1747 => x"06537573",
1748 => x"278d3888",
1749 => x"15085574",
1750 => x"782e0981",
1751 => x"06ea388c",
1752 => x"150880d5",
1753 => x"b40b8405",
1754 => x"08718c1a",
1755 => x"0c76881a",
1756 => x"0c788813",
1757 => x"0c788c18",
1758 => x"0c5d5879",
1759 => x"53807a24",
1760 => x"83e63872",
1761 => x"822c8171",
1762 => x"2b5c537a",
1763 => x"7c268198",
1764 => x"387b7b06",
1765 => x"537282f1",
1766 => x"3879fc06",
1767 => x"84055a7a",
1768 => x"10707d06",
1769 => x"545b7282",
1770 => x"e038841a",
1771 => x"5af13988",
1772 => x"178c1108",
1773 => x"58587678",
1774 => x"2e098106",
1775 => x"fcc23882",
1776 => x"1a5afdec",
1777 => x"39781779",
1778 => x"81078419",
1779 => x"0c7080d5",
1780 => x"c80c7080",
1781 => x"d5c40c80",
1782 => x"d5bc0b8c",
1783 => x"120c8c11",
1784 => x"0888120c",
1785 => x"74810784",
1786 => x"120c7411",
1787 => x"75710c51",
1788 => x"537d5188",
1789 => x"c63f8817",
1790 => x"54fcac39",
1791 => x"80d5b40b",
1792 => x"8405087a",
1793 => x"545c7980",
1794 => x"25fef838",
1795 => x"82da397a",
1796 => x"097c0670",
1797 => x"80d5b40b",
1798 => x"84050c5c",
1799 => x"7a105b7a",
1800 => x"7c268538",
1801 => x"7a85b838",
1802 => x"80d5b40b",
1803 => x"88050870",
1804 => x"841208fc",
1805 => x"06707c31",
1806 => x"7c72268f",
1807 => x"72250757",
1808 => x"575c5d55",
1809 => x"72802e80",
1810 => x"db38797a",
1811 => x"1680d5ac",
1812 => x"081b9011",
1813 => x"5a55575b",
1814 => x"80d5a808",
1815 => x"ff2e8838",
1816 => x"a08f13e0",
1817 => x"80065776",
1818 => x"527d5187",
1819 => x"cf3fb008",
1820 => x"54b008ff",
1821 => x"2e9038b0",
1822 => x"08762782",
1823 => x"99387480",
1824 => x"d5b42e82",
1825 => x"913880d5",
1826 => x"b40b8805",
1827 => x"08558415",
1828 => x"08fc0670",
1829 => x"7a317a72",
1830 => x"268f7225",
1831 => x"07525553",
1832 => x"7283e638",
1833 => x"74798107",
1834 => x"84170c79",
1835 => x"167080d5",
1836 => x"b40b8805",
1837 => x"0c758107",
1838 => x"84120c54",
1839 => x"7e525786",
1840 => x"fa3f8817",
1841 => x"54fae039",
1842 => x"75832a70",
1843 => x"54548074",
1844 => x"24819b38",
1845 => x"72822c81",
1846 => x"712b80d5",
1847 => x"b8080770",
1848 => x"80d5b40b",
1849 => x"84050c75",
1850 => x"10101080",
1851 => x"d5b40588",
1852 => x"1108585a",
1853 => x"5d53778c",
1854 => x"180c7488",
1855 => x"180c7688",
1856 => x"190c768c",
1857 => x"160cfcf3",
1858 => x"39797a10",
1859 => x"101080d5",
1860 => x"b4057057",
1861 => x"595d8c15",
1862 => x"08577675",
1863 => x"2ea33884",
1864 => x"1708fc06",
1865 => x"707a3155",
1866 => x"56738f24",
1867 => x"83ca3873",
1868 => x"80258481",
1869 => x"388c1708",
1870 => x"5776752e",
1871 => x"098106df",
1872 => x"38881581",
1873 => x"1b708306",
1874 => x"555b5572",
1875 => x"c9387c83",
1876 => x"06537280",
1877 => x"2efdb838",
1878 => x"ff1df819",
1879 => x"595d8818",
1880 => x"08782eea",
1881 => x"38fdb539",
1882 => x"831a53fc",
1883 => x"96398314",
1884 => x"70822c81",
1885 => x"712b80d5",
1886 => x"b8080770",
1887 => x"80d5b40b",
1888 => x"84050c76",
1889 => x"10101080",
1890 => x"d5b40588",
1891 => x"1108595b",
1892 => x"5e5153fe",
1893 => x"e13980d4",
1894 => x"f8081758",
1895 => x"b008762e",
1896 => x"818d3880",
1897 => x"d5a808ff",
1898 => x"2e83ec38",
1899 => x"73763118",
1900 => x"80d4f80c",
1901 => x"73870670",
1902 => x"57537280",
1903 => x"2e883888",
1904 => x"73317015",
1905 => x"55567614",
1906 => x"9fff06a0",
1907 => x"80713117",
1908 => x"70547f53",
1909 => x"575384e4",
1910 => x"3fb00853",
1911 => x"b008ff2e",
1912 => x"81a03880",
1913 => x"d4f80816",
1914 => x"7080d4f8",
1915 => x"0c747580",
1916 => x"d5b40b88",
1917 => x"050c7476",
1918 => x"31187081",
1919 => x"07515556",
1920 => x"587b80d5",
1921 => x"b42e839c",
1922 => x"38798f26",
1923 => x"82cb3881",
1924 => x"0b84150c",
1925 => x"841508fc",
1926 => x"06707a31",
1927 => x"7a72268f",
1928 => x"72250752",
1929 => x"55537280",
1930 => x"2efcf938",
1931 => x"80db39b0",
1932 => x"089fff06",
1933 => x"5372feeb",
1934 => x"387780d4",
1935 => x"f80c80d5",
1936 => x"b40b8805",
1937 => x"087b1881",
1938 => x"0784120c",
1939 => x"5580d5a4",
1940 => x"08782786",
1941 => x"387780d5",
1942 => x"a40c80d5",
1943 => x"a0087827",
1944 => x"fcac3877",
1945 => x"80d5a00c",
1946 => x"841508fc",
1947 => x"06707a31",
1948 => x"7a72268f",
1949 => x"72250752",
1950 => x"55537280",
1951 => x"2efca538",
1952 => x"88398074",
1953 => x"5456fedb",
1954 => x"397d5183",
1955 => x"ae3f800b",
1956 => x"b00c8f3d",
1957 => x"0d047353",
1958 => x"807424a9",
1959 => x"3872822c",
1960 => x"81712b80",
1961 => x"d5b80807",
1962 => x"7080d5b4",
1963 => x"0b84050c",
1964 => x"5d53778c",
1965 => x"180c7488",
1966 => x"180c7688",
1967 => x"190c768c",
1968 => x"160cf9b7",
1969 => x"39831470",
1970 => x"822c8171",
1971 => x"2b80d5b8",
1972 => x"08077080",
1973 => x"d5b40b84",
1974 => x"050c5e51",
1975 => x"53d4397b",
1976 => x"7b065372",
1977 => x"fca33884",
1978 => x"1a7b105c",
1979 => x"5af139ff",
1980 => x"1a811151",
1981 => x"5af7b939",
1982 => x"78177981",
1983 => x"0784190c",
1984 => x"8c180888",
1985 => x"1908718c",
1986 => x"120c8812",
1987 => x"0c597080",
1988 => x"d5c80c70",
1989 => x"80d5c40c",
1990 => x"80d5bc0b",
1991 => x"8c120c8c",
1992 => x"11088812",
1993 => x"0c748107",
1994 => x"84120c74",
1995 => x"1175710c",
1996 => x"5153f9bd",
1997 => x"39751784",
1998 => x"11088107",
1999 => x"84120c53",
2000 => x"8c170888",
2001 => x"1808718c",
2002 => x"120c8812",
2003 => x"0c587d51",
2004 => x"81e93f88",
2005 => x"1754f5cf",
2006 => x"39728415",
2007 => x"0cf41af8",
2008 => x"0670841e",
2009 => x"08810607",
2010 => x"841e0c70",
2011 => x"1d545b85",
2012 => x"0b84140c",
2013 => x"850b8814",
2014 => x"0c8f7b27",
2015 => x"fdcf3888",
2016 => x"1c527d51",
2017 => x"ec9e3f80",
2018 => x"d5b40b88",
2019 => x"050880d4",
2020 => x"f8085955",
2021 => x"fdb73977",
2022 => x"80d4f80c",
2023 => x"7380d5a8",
2024 => x"0cfc9139",
2025 => x"7284150c",
2026 => x"fda339fc",
2027 => x"3d0d7679",
2028 => x"71028c05",
2029 => x"9f053357",
2030 => x"55535583",
2031 => x"72278a38",
2032 => x"74830651",
2033 => x"70802ea2",
2034 => x"38ff1252",
2035 => x"71ff2e93",
2036 => x"38737370",
2037 => x"81055534",
2038 => x"ff125271",
2039 => x"ff2e0981",
2040 => x"06ef3874",
2041 => x"b00c863d",
2042 => x"0d047474",
2043 => x"882b7507",
2044 => x"7071902b",
2045 => x"07515451",
2046 => x"8f7227a5",
2047 => x"38727170",
2048 => x"8405530c",
2049 => x"72717084",
2050 => x"05530c72",
2051 => x"71708405",
2052 => x"530c7271",
2053 => x"70840553",
2054 => x"0cf01252",
2055 => x"718f26dd",
2056 => x"38837227",
2057 => x"90387271",
2058 => x"70840553",
2059 => x"0cfc1252",
2060 => x"718326f2",
2061 => x"387053ff",
2062 => x"90390404",
2063 => x"fd3d0d80",
2064 => x"0b80ddf4",
2065 => x"0c765184",
2066 => x"ee3fb008",
2067 => x"53b008ff",
2068 => x"2e883872",
2069 => x"b00c853d",
2070 => x"0d0480dd",
2071 => x"f4085473",
2072 => x"802ef038",
2073 => x"7574710c",
2074 => x"5272b00c",
2075 => x"853d0d04",
2076 => x"f93d0d79",
2077 => x"7c557b54",
2078 => x"8e112270",
2079 => x"902b7090",
2080 => x"2c555780",
2081 => x"cdf80853",
2082 => x"585683f3",
2083 => x"3fb00857",
2084 => x"800bb008",
2085 => x"24933880",
2086 => x"d01608b0",
2087 => x"080580d0",
2088 => x"170c76b0",
2089 => x"0c893d0d",
2090 => x"048c1622",
2091 => x"83dfff06",
2092 => x"55748c17",
2093 => x"2376b00c",
2094 => x"893d0d04",
2095 => x"fa3d0d78",
2096 => x"8c112270",
2097 => x"882a7081",
2098 => x"06515758",
2099 => x"5674a938",
2100 => x"8c162283",
2101 => x"dfff0655",
2102 => x"748c1723",
2103 => x"7a547953",
2104 => x"8e162270",
2105 => x"902b7090",
2106 => x"2c545680",
2107 => x"cdf80852",
2108 => x"5681b23f",
2109 => x"883d0d04",
2110 => x"82548053",
2111 => x"8e162270",
2112 => x"902b7090",
2113 => x"2c545680",
2114 => x"cdf80852",
2115 => x"5782b83f",
2116 => x"8c162283",
2117 => x"dfff0655",
2118 => x"748c1723",
2119 => x"7a547953",
2120 => x"8e162270",
2121 => x"902b7090",
2122 => x"2c545680",
2123 => x"cdf80852",
2124 => x"5680f23f",
2125 => x"883d0d04",
2126 => x"f93d0d79",
2127 => x"7c557b54",
2128 => x"8e112270",
2129 => x"902b7090",
2130 => x"2c555780",
2131 => x"cdf80853",
2132 => x"585681f3",
2133 => x"3fb00857",
2134 => x"b008ff2e",
2135 => x"99388c16",
2136 => x"22a08007",
2137 => x"55748c17",
2138 => x"23b00880",
2139 => x"d0170c76",
2140 => x"b00c893d",
2141 => x"0d048c16",
2142 => x"2283dfff",
2143 => x"0655748c",
2144 => x"172376b0",
2145 => x"0c893d0d",
2146 => x"04fe3d0d",
2147 => x"748e1122",
2148 => x"70902b70",
2149 => x"902c5551",
2150 => x"515380cd",
2151 => x"f80851bd",
2152 => x"3f843d0d",
2153 => x"04fb3d0d",
2154 => x"800b80dd",
2155 => x"f40c7a53",
2156 => x"79527851",
2157 => x"82fc3fb0",
2158 => x"0855b008",
2159 => x"ff2e8838",
2160 => x"74b00c87",
2161 => x"3d0d0480",
2162 => x"ddf40856",
2163 => x"75802ef0",
2164 => x"38777671",
2165 => x"0c5474b0",
2166 => x"0c873d0d",
2167 => x"04fd3d0d",
2168 => x"800b80dd",
2169 => x"f40c7651",
2170 => x"84c63fb0",
2171 => x"0853b008",
2172 => x"ff2e8838",
2173 => x"72b00c85",
2174 => x"3d0d0480",
2175 => x"ddf40854",
2176 => x"73802ef0",
2177 => x"38757471",
2178 => x"0c5272b0",
2179 => x"0c853d0d",
2180 => x"04fc3d0d",
2181 => x"800b80dd",
2182 => x"f40c7852",
2183 => x"775186ae",
2184 => x"3fb00854",
2185 => x"b008ff2e",
2186 => x"883873b0",
2187 => x"0c863d0d",
2188 => x"0480ddf4",
2189 => x"08557480",
2190 => x"2ef03876",
2191 => x"75710c53",
2192 => x"73b00c86",
2193 => x"3d0d04fb",
2194 => x"3d0d800b",
2195 => x"80ddf40c",
2196 => x"7a537952",
2197 => x"7851848a",
2198 => x"3fb00855",
2199 => x"b008ff2e",
2200 => x"883874b0",
2201 => x"0c873d0d",
2202 => x"0480ddf4",
2203 => x"08567580",
2204 => x"2ef03877",
2205 => x"76710c54",
2206 => x"74b00c87",
2207 => x"3d0d04fb",
2208 => x"3d0d800b",
2209 => x"80ddf40c",
2210 => x"7a537952",
2211 => x"78518296",
2212 => x"3fb00855",
2213 => x"b008ff2e",
2214 => x"883874b0",
2215 => x"0c873d0d",
2216 => x"0480ddf4",
2217 => x"08567580",
2218 => x"2ef03877",
2219 => x"76710c54",
2220 => x"74b00c87",
2221 => x"3d0d04fe",
2222 => x"3d0d80dd",
2223 => x"e4085170",
2224 => x"8a3880dd",
2225 => x"f87080dd",
2226 => x"e40c5170",
2227 => x"75125252",
2228 => x"ff537087",
2229 => x"fb808026",
2230 => x"88387080",
2231 => x"dde40c71",
2232 => x"5372b00c",
2233 => x"843d0d04",
2234 => x"fd3d0d80",
2235 => x"0b80cdec",
2236 => x"08545472",
2237 => x"812e9b38",
2238 => x"7380dde8",
2239 => x"0cc3e83f",
2240 => x"c1fe3f80",
2241 => x"ddbc5281",
2242 => x"51c5ac3f",
2243 => x"b0085185",
2244 => x"bd3f7280",
2245 => x"dde80cc3",
2246 => x"ce3fc1e4",
2247 => x"3f80ddbc",
2248 => x"528151c5",
2249 => x"923fb008",
2250 => x"5185a33f",
2251 => x"00ff3900",
2252 => x"ff39f53d",
2253 => x"0d7e6080",
2254 => x"dde80870",
2255 => x"5b585b5b",
2256 => x"7580c238",
2257 => x"777a25a1",
2258 => x"38771b70",
2259 => x"337081ff",
2260 => x"06585859",
2261 => x"758a2e98",
2262 => x"387681ff",
2263 => x"0651c2e6",
2264 => x"3f811858",
2265 => x"797824e1",
2266 => x"3879b00c",
2267 => x"8d3d0d04",
2268 => x"8d51c2d2",
2269 => x"3f783370",
2270 => x"81ff0652",
2271 => x"57c2c73f",
2272 => x"811858e0",
2273 => x"3979557a",
2274 => x"547d5385",
2275 => x"528d3dfc",
2276 => x"0551c1ae",
2277 => x"3fb00856",
2278 => x"84ad3f7b",
2279 => x"b0080c75",
2280 => x"b00c8d3d",
2281 => x"0d04f63d",
2282 => x"0d7d7f80",
2283 => x"dde80870",
2284 => x"5b585a5a",
2285 => x"7580c138",
2286 => x"777925b3",
2287 => x"38c1e23f",
2288 => x"b00881ff",
2289 => x"06708d32",
2290 => x"7030709f",
2291 => x"2a515157",
2292 => x"57768a2e",
2293 => x"80c33875",
2294 => x"802ebe38",
2295 => x"771a5676",
2296 => x"76347651",
2297 => x"c1e03f81",
2298 => x"18587878",
2299 => x"24cf3877",
2300 => x"5675b00c",
2301 => x"8c3d0d04",
2302 => x"78557954",
2303 => x"7c538452",
2304 => x"8c3dfc05",
2305 => x"51c0bb3f",
2306 => x"b0085683",
2307 => x"ba3f7ab0",
2308 => x"080c75b0",
2309 => x"0c8c3d0d",
2310 => x"04771a56",
2311 => x"8a763481",
2312 => x"18588d51",
2313 => x"c1a03f8a",
2314 => x"51c19b3f",
2315 => x"7756c239",
2316 => x"fb3d0d80",
2317 => x"dde80870",
2318 => x"56547388",
2319 => x"3874b00c",
2320 => x"873d0d04",
2321 => x"77538352",
2322 => x"873dfc05",
2323 => x"51ffbff2",
2324 => x"3fb00854",
2325 => x"82f13f75",
2326 => x"b0080c73",
2327 => x"b00c873d",
2328 => x"0d04fa3d",
2329 => x"0d80dde8",
2330 => x"08802ea3",
2331 => x"387a5579",
2332 => x"54785386",
2333 => x"52883dfc",
2334 => x"0551ffbf",
2335 => x"c53fb008",
2336 => x"5682c43f",
2337 => x"76b0080c",
2338 => x"75b00c88",
2339 => x"3d0d0482",
2340 => x"b63f9d0b",
2341 => x"b0080cff",
2342 => x"0bb00c88",
2343 => x"3d0d04fb",
2344 => x"3d0d7779",
2345 => x"56568070",
2346 => x"54547375",
2347 => x"259f3874",
2348 => x"101010f8",
2349 => x"05527216",
2350 => x"70337074",
2351 => x"2b760781",
2352 => x"16f81656",
2353 => x"56565151",
2354 => x"747324ea",
2355 => x"3873b00c",
2356 => x"873d0d04",
2357 => x"fc3d0d76",
2358 => x"785555bc",
2359 => x"53805273",
2360 => x"51f5c83f",
2361 => x"84527451",
2362 => x"ffb53fb0",
2363 => x"08742384",
2364 => x"52841551",
2365 => x"ffa93fb0",
2366 => x"08821523",
2367 => x"84528815",
2368 => x"51ff9c3f",
2369 => x"b0088415",
2370 => x"0c84528c",
2371 => x"1551ff8f",
2372 => x"3fb00888",
2373 => x"15238452",
2374 => x"901551ff",
2375 => x"823fb008",
2376 => x"8a152384",
2377 => x"52941551",
2378 => x"fef53fb0",
2379 => x"088c1523",
2380 => x"84529815",
2381 => x"51fee83f",
2382 => x"b0088e15",
2383 => x"2388529c",
2384 => x"1551fedb",
2385 => x"3fb00890",
2386 => x"150c863d",
2387 => x"0d04e93d",
2388 => x"0d6a80dd",
2389 => x"e8085757",
2390 => x"75933880",
2391 => x"c0800b84",
2392 => x"180c75ac",
2393 => x"180c75b0",
2394 => x"0c993d0d",
2395 => x"04893d70",
2396 => x"556a5455",
2397 => x"8a52993d",
2398 => x"ffbc0551",
2399 => x"ffbdc33f",
2400 => x"b0087753",
2401 => x"755256fe",
2402 => x"cb3fbc3f",
2403 => x"77b0080c",
2404 => x"75b00c99",
2405 => x"3d0d04fc",
2406 => x"3d0d8154",
2407 => x"80dde808",
2408 => x"883873b0",
2409 => x"0c863d0d",
2410 => x"04765397",
2411 => x"b952863d",
2412 => x"fc0551ff",
2413 => x"bd8c3fb0",
2414 => x"08548c3f",
2415 => x"74b0080c",
2416 => x"73b00c86",
2417 => x"3d0d0480",
2418 => x"cdf808b0",
2419 => x"0c04f73d",
2420 => x"0d7b80cd",
2421 => x"f80882c8",
2422 => x"11085a54",
2423 => x"5a77802e",
2424 => x"80da3881",
2425 => x"88188419",
2426 => x"08ff0581",
2427 => x"712b5955",
2428 => x"59807424",
2429 => x"80ea3880",
2430 => x"7424b538",
2431 => x"73822b78",
2432 => x"11880556",
2433 => x"56818019",
2434 => x"08770653",
2435 => x"72802eb6",
2436 => x"38781670",
2437 => x"08535379",
2438 => x"51740853",
2439 => x"722dff14",
2440 => x"fc17fc17",
2441 => x"79812c5a",
2442 => x"57575473",
2443 => x"8025d638",
2444 => x"77085877",
2445 => x"ffad3880",
2446 => x"cdf80853",
2447 => x"bc1308a5",
2448 => x"387951f9",
2449 => x"e73f7408",
2450 => x"53722dff",
2451 => x"14fc17fc",
2452 => x"1779812c",
2453 => x"5a575754",
2454 => x"738025ff",
2455 => x"a838d139",
2456 => x"8057ff93",
2457 => x"397251bc",
2458 => x"13085372",
2459 => x"2d7951f9",
2460 => x"bb3fff3d",
2461 => x"0d80ddc4",
2462 => x"0bfc0570",
2463 => x"08525270",
2464 => x"ff2e9138",
2465 => x"702dfc12",
2466 => x"70085252",
2467 => x"70ff2e09",
2468 => x"8106f138",
2469 => x"833d0d04",
2470 => x"04ffbdb6",
2471 => x"3f040000",
2472 => x"00ffffff",
2473 => x"ff00ffff",
2474 => x"ffff00ff",
2475 => x"ffffff00",
2476 => x"00000040",
2477 => x"48656c6c",
2478 => x"6f20776f",
2479 => x"726c6420",
2480 => x"310a0000",
2481 => x"48656c6c",
2482 => x"6f20776f",
2483 => x"726c6420",
2484 => x"320a0000",
2485 => x"0a000000",
2486 => x"43000000",
2487 => x"64756d6d",
2488 => x"792e6578",
2489 => x"65000000",
2490 => x"00000000",
2491 => x"00000000",
2492 => x"00000000",
2493 => x"00002ecc",
2494 => x"000026fc",
2495 => x"00000000",
2496 => x"00002964",
2497 => x"000029c0",
2498 => x"00002a1c",
2499 => x"00000000",
2500 => x"00000000",
2501 => x"00000000",
2502 => x"00000000",
2503 => x"00000000",
2504 => x"00000000",
2505 => x"00000000",
2506 => x"00000000",
2507 => x"00000000",
2508 => x"000026d8",
2509 => x"00000000",
2510 => x"00000000",
2511 => x"00000000",
2512 => x"00000000",
2513 => x"00000000",
2514 => x"00000000",
2515 => x"00000000",
2516 => x"00000000",
2517 => x"00000000",
2518 => x"00000000",
2519 => x"00000000",
2520 => x"00000000",
2521 => x"00000000",
2522 => x"00000000",
2523 => x"00000000",
2524 => x"00000000",
2525 => x"00000000",
2526 => x"00000000",
2527 => x"00000000",
2528 => x"00000000",
2529 => x"00000000",
2530 => x"00000000",
2531 => x"00000000",
2532 => x"00000000",
2533 => x"00000000",
2534 => x"00000000",
2535 => x"00000000",
2536 => x"00000000",
2537 => x"00000001",
2538 => x"330eabcd",
2539 => x"1234e66d",
2540 => x"deec0005",
2541 => x"000b0000",
2542 => x"00000000",
2543 => x"00000000",
2544 => x"00000000",
2545 => x"00000000",
2546 => x"00000000",
2547 => x"00000000",
2548 => x"00000000",
2549 => x"00000000",
2550 => x"00000000",
2551 => x"00000000",
2552 => x"00000000",
2553 => x"00000000",
2554 => x"00000000",
2555 => x"00000000",
2556 => x"00000000",
2557 => x"00000000",
2558 => x"00000000",
2559 => x"00000000",
2560 => x"00000000",
2561 => x"00000000",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"00000000",
2568 => x"00000000",
2569 => x"00000000",
2570 => x"00000000",
2571 => x"00000000",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000000",
2586 => x"00000000",
2587 => x"00000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000000",
2597 => x"00000000",
2598 => x"00000000",
2599 => x"00000000",
2600 => x"00000000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"ffffffff",
2731 => x"00000000",
2732 => x"00020000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00002ab4",
2736 => x"00002ab4",
2737 => x"00002abc",
2738 => x"00002abc",
2739 => x"00002ac4",
2740 => x"00002ac4",
2741 => x"00002acc",
2742 => x"00002acc",
2743 => x"00002ad4",
2744 => x"00002ad4",
2745 => x"00002adc",
2746 => x"00002adc",
2747 => x"00002ae4",
2748 => x"00002ae4",
2749 => x"00002aec",
2750 => x"00002aec",
2751 => x"00002af4",
2752 => x"00002af4",
2753 => x"00002afc",
2754 => x"00002afc",
2755 => x"00002b04",
2756 => x"00002b04",
2757 => x"00002b0c",
2758 => x"00002b0c",
2759 => x"00002b14",
2760 => x"00002b14",
2761 => x"00002b1c",
2762 => x"00002b1c",
2763 => x"00002b24",
2764 => x"00002b24",
2765 => x"00002b2c",
2766 => x"00002b2c",
2767 => x"00002b34",
2768 => x"00002b34",
2769 => x"00002b3c",
2770 => x"00002b3c",
2771 => x"00002b44",
2772 => x"00002b44",
2773 => x"00002b4c",
2774 => x"00002b4c",
2775 => x"00002b54",
2776 => x"00002b54",
2777 => x"00002b5c",
2778 => x"00002b5c",
2779 => x"00002b64",
2780 => x"00002b64",
2781 => x"00002b6c",
2782 => x"00002b6c",
2783 => x"00002b74",
2784 => x"00002b74",
2785 => x"00002b7c",
2786 => x"00002b7c",
2787 => x"00002b84",
2788 => x"00002b84",
2789 => x"00002b8c",
2790 => x"00002b8c",
2791 => x"00002b94",
2792 => x"00002b94",
2793 => x"00002b9c",
2794 => x"00002b9c",
2795 => x"00002ba4",
2796 => x"00002ba4",
2797 => x"00002bac",
2798 => x"00002bac",
2799 => x"00002bb4",
2800 => x"00002bb4",
2801 => x"00002bbc",
2802 => x"00002bbc",
2803 => x"00002bc4",
2804 => x"00002bc4",
2805 => x"00002bcc",
2806 => x"00002bcc",
2807 => x"00002bd4",
2808 => x"00002bd4",
2809 => x"00002bdc",
2810 => x"00002bdc",
2811 => x"00002be4",
2812 => x"00002be4",
2813 => x"00002bec",
2814 => x"00002bec",
2815 => x"00002bf4",
2816 => x"00002bf4",
2817 => x"00002bfc",
2818 => x"00002bfc",
2819 => x"00002c04",
2820 => x"00002c04",
2821 => x"00002c0c",
2822 => x"00002c0c",
2823 => x"00002c14",
2824 => x"00002c14",
2825 => x"00002c1c",
2826 => x"00002c1c",
2827 => x"00002c24",
2828 => x"00002c24",
2829 => x"00002c2c",
2830 => x"00002c2c",
2831 => x"00002c34",
2832 => x"00002c34",
2833 => x"00002c3c",
2834 => x"00002c3c",
2835 => x"00002c44",
2836 => x"00002c44",
2837 => x"00002c4c",
2838 => x"00002c4c",
2839 => x"00002c54",
2840 => x"00002c54",
2841 => x"00002c5c",
2842 => x"00002c5c",
2843 => x"00002c64",
2844 => x"00002c64",
2845 => x"00002c6c",
2846 => x"00002c6c",
2847 => x"00002c74",
2848 => x"00002c74",
2849 => x"00002c7c",
2850 => x"00002c7c",
2851 => x"00002c84",
2852 => x"00002c84",
2853 => x"00002c8c",
2854 => x"00002c8c",
2855 => x"00002c94",
2856 => x"00002c94",
2857 => x"00002c9c",
2858 => x"00002c9c",
2859 => x"00002ca4",
2860 => x"00002ca4",
2861 => x"00002cac",
2862 => x"00002cac",
2863 => x"00002cb4",
2864 => x"00002cb4",
2865 => x"00002cbc",
2866 => x"00002cbc",
2867 => x"00002cc4",
2868 => x"00002cc4",
2869 => x"00002ccc",
2870 => x"00002ccc",
2871 => x"00002cd4",
2872 => x"00002cd4",
2873 => x"00002cdc",
2874 => x"00002cdc",
2875 => x"00002ce4",
2876 => x"00002ce4",
2877 => x"00002cec",
2878 => x"00002cec",
2879 => x"00002cf4",
2880 => x"00002cf4",
2881 => x"00002cfc",
2882 => x"00002cfc",
2883 => x"00002d04",
2884 => x"00002d04",
2885 => x"00002d0c",
2886 => x"00002d0c",
2887 => x"00002d14",
2888 => x"00002d14",
2889 => x"00002d1c",
2890 => x"00002d1c",
2891 => x"00002d24",
2892 => x"00002d24",
2893 => x"00002d2c",
2894 => x"00002d2c",
2895 => x"00002d34",
2896 => x"00002d34",
2897 => x"00002d3c",
2898 => x"00002d3c",
2899 => x"00002d44",
2900 => x"00002d44",
2901 => x"00002d4c",
2902 => x"00002d4c",
2903 => x"00002d54",
2904 => x"00002d54",
2905 => x"00002d5c",
2906 => x"00002d5c",
2907 => x"00002d64",
2908 => x"00002d64",
2909 => x"00002d6c",
2910 => x"00002d6c",
2911 => x"00002d74",
2912 => x"00002d74",
2913 => x"00002d7c",
2914 => x"00002d7c",
2915 => x"00002d84",
2916 => x"00002d84",
2917 => x"00002d8c",
2918 => x"00002d8c",
2919 => x"00002d94",
2920 => x"00002d94",
2921 => x"00002d9c",
2922 => x"00002d9c",
2923 => x"00002da4",
2924 => x"00002da4",
2925 => x"00002dac",
2926 => x"00002dac",
2927 => x"00002db4",
2928 => x"00002db4",
2929 => x"00002dbc",
2930 => x"00002dbc",
2931 => x"00002dc4",
2932 => x"00002dc4",
2933 => x"00002dcc",
2934 => x"00002dcc",
2935 => x"00002dd4",
2936 => x"00002dd4",
2937 => x"00002ddc",
2938 => x"00002ddc",
2939 => x"00002de4",
2940 => x"00002de4",
2941 => x"00002dec",
2942 => x"00002dec",
2943 => x"00002df4",
2944 => x"00002df4",
2945 => x"00002dfc",
2946 => x"00002dfc",
2947 => x"00002e04",
2948 => x"00002e04",
2949 => x"00002e0c",
2950 => x"00002e0c",
2951 => x"00002e14",
2952 => x"00002e14",
2953 => x"00002e1c",
2954 => x"00002e1c",
2955 => x"00002e24",
2956 => x"00002e24",
2957 => x"00002e2c",
2958 => x"00002e2c",
2959 => x"00002e34",
2960 => x"00002e34",
2961 => x"00002e3c",
2962 => x"00002e3c",
2963 => x"00002e44",
2964 => x"00002e44",
2965 => x"00002e4c",
2966 => x"00002e4c",
2967 => x"00002e54",
2968 => x"00002e54",
2969 => x"00002e5c",
2970 => x"00002e5c",
2971 => x"00002e64",
2972 => x"00002e64",
2973 => x"00002e6c",
2974 => x"00002e6c",
2975 => x"00002e74",
2976 => x"00002e74",
2977 => x"00002e7c",
2978 => x"00002e7c",
2979 => x"00002e84",
2980 => x"00002e84",
2981 => x"00002e8c",
2982 => x"00002e8c",
2983 => x"00002e94",
2984 => x"00002e94",
2985 => x"00002e9c",
2986 => x"00002e9c",
2987 => x"00002ea4",
2988 => x"00002ea4",
2989 => x"00002eac",
2990 => x"00002eac",
2991 => x"000026dc",
2992 => x"ffffffff",
2993 => x"00000000",
2994 => x"ffffffff",
2995 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

