------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80d1b80c",
3 => x"3a0b0b80",
4 => x"c9ab0400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d0",
162 => x"ec738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d1b40c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c8b93f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"90db2d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8fa92d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80e1a4",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80e1",
307 => x"a4085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480d1",
314 => x"b408802e",
315 => x"a43880d1",
316 => x"b808822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80e1a40c",
320 => x"82a0800b",
321 => x"80e1a80c",
322 => x"8290800b",
323 => x"80e1ac0c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80e1a4",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"e1a80cf8",
330 => x"80808480",
331 => x"0b80e1ac",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80e1",
335 => x"a40c80c0",
336 => x"a880940b",
337 => x"80e1a80c",
338 => x"80d0fc0b",
339 => x"80e1ac0c",
340 => x"04ff3d0d",
341 => x"80e1b033",
342 => x"5170a738",
343 => x"80d1c008",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"d1c00c70",
348 => x"2d80d1c0",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80e1",
352 => x"b034833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80e1a008",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"e1a0510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404803d",
366 => x"0d80e1bc",
367 => x"08811180",
368 => x"e1bc0c51",
369 => x"823d0d04",
370 => x"f73d0d7b",
371 => x"54870b89",
372 => x"3d80d1c4",
373 => x"08585855",
374 => x"7417748f",
375 => x"06175353",
376 => x"71337334",
377 => x"73842aff",
378 => x"16565474",
379 => x"8025e938",
380 => x"800b8b3d",
381 => x"34765189",
382 => x"853f8b3d",
383 => x"0d04e13d",
384 => x"0d80e1bc",
385 => x"089f3d9d",
386 => x"3d9b3d99",
387 => x"3d973d95",
388 => x"3d8c8080",
389 => x"088c8084",
390 => x"088e8080",
391 => x"0880d194",
392 => x"5b415f57",
393 => x"5f5f5f5f",
394 => x"5f5f5288",
395 => x"d13f7154",
396 => x"870b80d1",
397 => x"c4085755",
398 => x"741e748f",
399 => x"06175353",
400 => x"71337334",
401 => x"73842aff",
402 => x"16565474",
403 => x"8025e938",
404 => x"800ba13d",
405 => x"347d5188",
406 => x"a53f80d1",
407 => x"9851889e",
408 => x"3f765487",
409 => x"0b80d1c4",
410 => x"08575574",
411 => x"1d748f06",
412 => x"17545772",
413 => x"33773473",
414 => x"842aff16",
415 => x"56547480",
416 => x"25e93880",
417 => x"0b9e3d34",
418 => x"7c5187f2",
419 => x"3f80d19c",
420 => x"5187eb3f",
421 => x"7754870b",
422 => x"80d1c408",
423 => x"5755741c",
424 => x"748f0617",
425 => x"53587133",
426 => x"78347384",
427 => x"2aff1656",
428 => x"54748025",
429 => x"e938800b",
430 => x"9b3d347b",
431 => x"5187bf3f",
432 => x"f8bb9586",
433 => x"a10b8c80",
434 => x"800c8191",
435 => x"d1acf80b",
436 => x"8c80840c",
437 => x"f9d5f3bd",
438 => x"f00b8e80",
439 => x"800c8c80",
440 => x"80088c80",
441 => x"84088e80",
442 => x"800880d1",
443 => x"94545a58",
444 => x"55878b3f",
445 => x"7454870b",
446 => x"80d1c408",
447 => x"5755741b",
448 => x"748f0617",
449 => x"53537133",
450 => x"73347384",
451 => x"2aff1656",
452 => x"54748025",
453 => x"e938800b",
454 => x"983d347a",
455 => x"5186df3f",
456 => x"80d19851",
457 => x"86d83f76",
458 => x"54870b80",
459 => x"d1c40857",
460 => x"55741a74",
461 => x"8f061754",
462 => x"57723377",
463 => x"3473842a",
464 => x"ff165654",
465 => x"748025e9",
466 => x"38800b95",
467 => x"3d347951",
468 => x"86ac3f80",
469 => x"d19c5186",
470 => x"a53f7754",
471 => x"870b80d1",
472 => x"c4085755",
473 => x"7419748f",
474 => x"06175358",
475 => x"71337834",
476 => x"73842aff",
477 => x"16565474",
478 => x"8025e938",
479 => x"800b923d",
480 => x"34785185",
481 => x"f93f8c80",
482 => x"80088c80",
483 => x"84088e80",
484 => x"800880d1",
485 => x"94545a58",
486 => x"5285e33f",
487 => x"7154870b",
488 => x"80d1c408",
489 => x"5755fd90",
490 => x"39bc0802",
491 => x"bc0cf93d",
492 => x"0d800bbc",
493 => x"08fc050c",
494 => x"bc088805",
495 => x"088025ab",
496 => x"38bc0888",
497 => x"050830bc",
498 => x"0888050c",
499 => x"800bbc08",
500 => x"f4050cbc",
501 => x"08fc0508",
502 => x"8838810b",
503 => x"bc08f405",
504 => x"0cbc08f4",
505 => x"0508bc08",
506 => x"fc050cbc",
507 => x"088c0508",
508 => x"8025ab38",
509 => x"bc088c05",
510 => x"0830bc08",
511 => x"8c050c80",
512 => x"0bbc08f0",
513 => x"050cbc08",
514 => x"fc050888",
515 => x"38810bbc",
516 => x"08f0050c",
517 => x"bc08f005",
518 => x"08bc08fc",
519 => x"050c8053",
520 => x"bc088c05",
521 => x"0852bc08",
522 => x"88050851",
523 => x"81a73fb0",
524 => x"0870bc08",
525 => x"f8050c54",
526 => x"bc08fc05",
527 => x"08802e8c",
528 => x"38bc08f8",
529 => x"050830bc",
530 => x"08f8050c",
531 => x"bc08f805",
532 => x"0870b00c",
533 => x"54893d0d",
534 => x"bc0c04bc",
535 => x"0802bc0c",
536 => x"fb3d0d80",
537 => x"0bbc08fc",
538 => x"050cbc08",
539 => x"88050880",
540 => x"259338bc",
541 => x"08880508",
542 => x"30bc0888",
543 => x"050c810b",
544 => x"bc08fc05",
545 => x"0cbc088c",
546 => x"05088025",
547 => x"8c38bc08",
548 => x"8c050830",
549 => x"bc088c05",
550 => x"0c8153bc",
551 => x"088c0508",
552 => x"52bc0888",
553 => x"050851ad",
554 => x"3fb00870",
555 => x"bc08f805",
556 => x"0c54bc08",
557 => x"fc050880",
558 => x"2e8c38bc",
559 => x"08f80508",
560 => x"30bc08f8",
561 => x"050cbc08",
562 => x"f8050870",
563 => x"b00c5487",
564 => x"3d0dbc0c",
565 => x"04bc0802",
566 => x"bc0cfd3d",
567 => x"0d810bbc",
568 => x"08fc050c",
569 => x"800bbc08",
570 => x"f8050cbc",
571 => x"088c0508",
572 => x"bc088805",
573 => x"0827ac38",
574 => x"bc08fc05",
575 => x"08802ea3",
576 => x"38800bbc",
577 => x"088c0508",
578 => x"249938bc",
579 => x"088c0508",
580 => x"10bc088c",
581 => x"050cbc08",
582 => x"fc050810",
583 => x"bc08fc05",
584 => x"0cc939bc",
585 => x"08fc0508",
586 => x"802e80c9",
587 => x"38bc088c",
588 => x"0508bc08",
589 => x"88050826",
590 => x"a138bc08",
591 => x"880508bc",
592 => x"088c0508",
593 => x"31bc0888",
594 => x"050cbc08",
595 => x"f80508bc",
596 => x"08fc0508",
597 => x"07bc08f8",
598 => x"050cbc08",
599 => x"fc050881",
600 => x"2abc08fc",
601 => x"050cbc08",
602 => x"8c050881",
603 => x"2abc088c",
604 => x"050cffaf",
605 => x"39bc0890",
606 => x"0508802e",
607 => x"8f38bc08",
608 => x"88050870",
609 => x"bc08f405",
610 => x"0c518d39",
611 => x"bc08f805",
612 => x"0870bc08",
613 => x"f4050c51",
614 => x"bc08f405",
615 => x"08b00c85",
616 => x"3d0dbc0c",
617 => x"04fc3d0d",
618 => x"7670797b",
619 => x"55555555",
620 => x"8f72278c",
621 => x"38727507",
622 => x"83065170",
623 => x"802ea738",
624 => x"ff125271",
625 => x"ff2e9838",
626 => x"72708105",
627 => x"54337470",
628 => x"81055634",
629 => x"ff125271",
630 => x"ff2e0981",
631 => x"06ea3874",
632 => x"b00c863d",
633 => x"0d047451",
634 => x"72708405",
635 => x"54087170",
636 => x"8405530c",
637 => x"72708405",
638 => x"54087170",
639 => x"8405530c",
640 => x"72708405",
641 => x"54087170",
642 => x"8405530c",
643 => x"72708405",
644 => x"54087170",
645 => x"8405530c",
646 => x"f0125271",
647 => x"8f26c938",
648 => x"83722795",
649 => x"38727084",
650 => x"05540871",
651 => x"70840553",
652 => x"0cfc1252",
653 => x"718326ed",
654 => x"387054ff",
655 => x"8339f73d",
656 => x"0d7c7052",
657 => x"5380c83f",
658 => x"7254b008",
659 => x"5580d1a0",
660 => x"568157b0",
661 => x"0881055a",
662 => x"8b3de411",
663 => x"59538259",
664 => x"f413527b",
665 => x"88110852",
666 => x"5381833f",
667 => x"b0083070",
668 => x"b008079f",
669 => x"2c8a07b0",
670 => x"0c538b3d",
671 => x"0d04ff3d",
672 => x"0d735280",
673 => x"d1c80851",
674 => x"ffb43f83",
675 => x"3d0d04fd",
676 => x"3d0d7570",
677 => x"71830653",
678 => x"555270b8",
679 => x"38717008",
680 => x"7009f7fb",
681 => x"fdff1206",
682 => x"70f88482",
683 => x"81800651",
684 => x"51525370",
685 => x"9d388413",
686 => x"70087009",
687 => x"f7fbfdff",
688 => x"120670f8",
689 => x"84828180",
690 => x"06515152",
691 => x"5370802e",
692 => x"e5387252",
693 => x"71335170",
694 => x"802e8a38",
695 => x"81127033",
696 => x"525270f8",
697 => x"38717431",
698 => x"b00c853d",
699 => x"0d04f23d",
700 => x"0d606288",
701 => x"11087057",
702 => x"575f5a74",
703 => x"802e818f",
704 => x"388c1a22",
705 => x"70832a81",
706 => x"32708106",
707 => x"51555873",
708 => x"8638901a",
709 => x"08913879",
710 => x"5190a13f",
711 => x"ff54b008",
712 => x"80ed388c",
713 => x"1a22587d",
714 => x"08578078",
715 => x"83ffff06",
716 => x"70812a70",
717 => x"81065156",
718 => x"57557375",
719 => x"2e80d738",
720 => x"74903876",
721 => x"08841808",
722 => x"88195956",
723 => x"5974802e",
724 => x"f2387454",
725 => x"88807527",
726 => x"84388880",
727 => x"54735378",
728 => x"529c1a08",
729 => x"51a41a08",
730 => x"54732d80",
731 => x"0bb00825",
732 => x"82e638b0",
733 => x"081975b0",
734 => x"08317f88",
735 => x"0508b008",
736 => x"31706188",
737 => x"050c5656",
738 => x"5973ffb4",
739 => x"38805473",
740 => x"b00c903d",
741 => x"0d047581",
742 => x"32708106",
743 => x"76415154",
744 => x"73802e81",
745 => x"c1387490",
746 => x"38760884",
747 => x"18088819",
748 => x"59565974",
749 => x"802ef238",
750 => x"881a0878",
751 => x"83ffff06",
752 => x"70892a70",
753 => x"81065156",
754 => x"59567380",
755 => x"2e82fa38",
756 => x"7575278d",
757 => x"3877872a",
758 => x"70810651",
759 => x"547382b5",
760 => x"38747627",
761 => x"83387456",
762 => x"75537852",
763 => x"79085185",
764 => x"823f881a",
765 => x"08763188",
766 => x"1b0c7908",
767 => x"167a0c74",
768 => x"56751975",
769 => x"77317f88",
770 => x"05087831",
771 => x"70618805",
772 => x"0c565659",
773 => x"73802efe",
774 => x"f4388c1a",
775 => x"2258ff86",
776 => x"39777854",
777 => x"79537b52",
778 => x"5684c83f",
779 => x"881a0878",
780 => x"31881b0c",
781 => x"7908187a",
782 => x"0c7c7631",
783 => x"5d7c8e38",
784 => x"79518fdb",
785 => x"3fb00881",
786 => x"8f38b008",
787 => x"5f751975",
788 => x"77317f88",
789 => x"05087831",
790 => x"70618805",
791 => x"0c565659",
792 => x"73802efe",
793 => x"a8387481",
794 => x"83387608",
795 => x"84180888",
796 => x"19595659",
797 => x"74802ef2",
798 => x"3874538a",
799 => x"52785182",
800 => x"d33fb008",
801 => x"79318105",
802 => x"5db00884",
803 => x"3881155d",
804 => x"815f7c58",
805 => x"747d2783",
806 => x"38745894",
807 => x"1a08881b",
808 => x"0811575c",
809 => x"807a085c",
810 => x"54901a08",
811 => x"7b278338",
812 => x"81547578",
813 => x"25843873",
814 => x"ba387b78",
815 => x"24fee238",
816 => x"7b537852",
817 => x"9c1a0851",
818 => x"a41a0854",
819 => x"732db008",
820 => x"56b00880",
821 => x"24fee238",
822 => x"8c1a2280",
823 => x"c0075473",
824 => x"8c1b23ff",
825 => x"5473b00c",
826 => x"903d0d04",
827 => x"7effa338",
828 => x"ff873975",
829 => x"5378527a",
830 => x"5182f83f",
831 => x"7908167a",
832 => x"0c79518e",
833 => x"9a3fb008",
834 => x"cf387c76",
835 => x"315d7cfe",
836 => x"bc38feac",
837 => x"39901a08",
838 => x"7a087131",
839 => x"76117056",
840 => x"5a575280",
841 => x"d1c80851",
842 => x"848c3fb0",
843 => x"08802eff",
844 => x"a738b008",
845 => x"901b0cb0",
846 => x"08167a0c",
847 => x"77941b0c",
848 => x"74881b0c",
849 => x"7456fd99",
850 => x"39790858",
851 => x"901a0878",
852 => x"27833881",
853 => x"54757527",
854 => x"843873b3",
855 => x"38941a08",
856 => x"56757526",
857 => x"80d33875",
858 => x"5378529c",
859 => x"1a0851a4",
860 => x"1a085473",
861 => x"2db00856",
862 => x"b0088024",
863 => x"fd83388c",
864 => x"1a2280c0",
865 => x"0754738c",
866 => x"1b23ff54",
867 => x"fed73975",
868 => x"53785277",
869 => x"5181dc3f",
870 => x"7908167a",
871 => x"0c79518c",
872 => x"fe3fb008",
873 => x"802efcd9",
874 => x"388c1a22",
875 => x"80c00754",
876 => x"738c1b23",
877 => x"ff54fead",
878 => x"39747554",
879 => x"79537852",
880 => x"5681b03f",
881 => x"881a0875",
882 => x"31881b0c",
883 => x"7908157a",
884 => x"0cfcae39",
885 => x"fa3d0d7a",
886 => x"79028805",
887 => x"a7053356",
888 => x"52538373",
889 => x"278a3870",
890 => x"83065271",
891 => x"802ea838",
892 => x"ff135372",
893 => x"ff2e9738",
894 => x"70335273",
895 => x"722e9138",
896 => x"8111ff14",
897 => x"545172ff",
898 => x"2e098106",
899 => x"eb388051",
900 => x"70b00c88",
901 => x"3d0d0470",
902 => x"72575583",
903 => x"51758280",
904 => x"2914ff12",
905 => x"52567080",
906 => x"25f33883",
907 => x"7327bf38",
908 => x"74087632",
909 => x"7009f7fb",
910 => x"fdff1206",
911 => x"70f88482",
912 => x"81800651",
913 => x"51517080",
914 => x"2e993874",
915 => x"51805270",
916 => x"33577377",
917 => x"2effb938",
918 => x"81118113",
919 => x"53518372",
920 => x"27ed38fc",
921 => x"13841656",
922 => x"53728326",
923 => x"c3387451",
924 => x"fefe39fa",
925 => x"3d0d787a",
926 => x"7c727272",
927 => x"57575759",
928 => x"56567476",
929 => x"27b23876",
930 => x"15517571",
931 => x"27aa3870",
932 => x"7717ff14",
933 => x"54555371",
934 => x"ff2e9638",
935 => x"ff14ff14",
936 => x"54547233",
937 => x"7434ff12",
938 => x"5271ff2e",
939 => x"098106ec",
940 => x"3875b00c",
941 => x"883d0d04",
942 => x"768f2697",
943 => x"38ff1252",
944 => x"71ff2eed",
945 => x"38727081",
946 => x"05543374",
947 => x"70810556",
948 => x"34eb3974",
949 => x"76078306",
950 => x"5170e238",
951 => x"75755451",
952 => x"72708405",
953 => x"54087170",
954 => x"8405530c",
955 => x"72708405",
956 => x"54087170",
957 => x"8405530c",
958 => x"72708405",
959 => x"54087170",
960 => x"8405530c",
961 => x"72708405",
962 => x"54087170",
963 => x"8405530c",
964 => x"f0125271",
965 => x"8f26c938",
966 => x"83722795",
967 => x"38727084",
968 => x"05540871",
969 => x"70840553",
970 => x"0cfc1252",
971 => x"718326ed",
972 => x"387054ff",
973 => x"8839ef3d",
974 => x"0d636567",
975 => x"405d427b",
976 => x"802e84fa",
977 => x"386151a5",
978 => x"b43ff81c",
979 => x"70841208",
980 => x"70fc0670",
981 => x"628b0570",
982 => x"f8064159",
983 => x"455b5c41",
984 => x"57967427",
985 => x"82c33880",
986 => x"7b247e7c",
987 => x"26075980",
988 => x"5478742e",
989 => x"09810682",
990 => x"a938777b",
991 => x"2581fc38",
992 => x"771780d9",
993 => x"840b8805",
994 => x"085e567c",
995 => x"762e84bd",
996 => x"38841608",
997 => x"70fe0617",
998 => x"84110881",
999 => x"06515555",
1000 => x"73828b38",
1001 => x"74fc0659",
1002 => x"7c762e84",
1003 => x"dd387719",
1004 => x"5f7e7b25",
1005 => x"81fd3879",
1006 => x"81065473",
1007 => x"82bf3876",
1008 => x"77083184",
1009 => x"1108fc06",
1010 => x"565a7580",
1011 => x"2e91387c",
1012 => x"762e84ea",
1013 => x"38741918",
1014 => x"59787b25",
1015 => x"84893879",
1016 => x"802e8299",
1017 => x"38771556",
1018 => x"7a762482",
1019 => x"90388c1a",
1020 => x"08881b08",
1021 => x"718c120c",
1022 => x"88120c55",
1023 => x"79765957",
1024 => x"881761fc",
1025 => x"05575975",
1026 => x"a42685ef",
1027 => x"387b7955",
1028 => x"55937627",
1029 => x"80c9387b",
1030 => x"7084055d",
1031 => x"087c5679",
1032 => x"0c747084",
1033 => x"0556088c",
1034 => x"180c9017",
1035 => x"549b7627",
1036 => x"ae387470",
1037 => x"84055608",
1038 => x"740c7470",
1039 => x"84055608",
1040 => x"94180c98",
1041 => x"1754a376",
1042 => x"27953874",
1043 => x"70840556",
1044 => x"08740c74",
1045 => x"70840556",
1046 => x"089c180c",
1047 => x"a0175474",
1048 => x"70840556",
1049 => x"08747084",
1050 => x"05560c74",
1051 => x"70840556",
1052 => x"08747084",
1053 => x"05560c74",
1054 => x"08740c77",
1055 => x"7b315675",
1056 => x"8f2680c9",
1057 => x"38841708",
1058 => x"81067807",
1059 => x"84180c77",
1060 => x"17841108",
1061 => x"81078412",
1062 => x"0c546151",
1063 => x"a2e03f88",
1064 => x"175473b0",
1065 => x"0c933d0d",
1066 => x"04905bfd",
1067 => x"ba397856",
1068 => x"fe85398c",
1069 => x"16088817",
1070 => x"08718c12",
1071 => x"0c88120c",
1072 => x"557e707c",
1073 => x"3157588f",
1074 => x"7627ffb9",
1075 => x"387a1784",
1076 => x"18088106",
1077 => x"7c078419",
1078 => x"0c768107",
1079 => x"84120c76",
1080 => x"11841108",
1081 => x"81078412",
1082 => x"0c558805",
1083 => x"5261518c",
1084 => x"f63f6151",
1085 => x"a2883f88",
1086 => x"1754ffa6",
1087 => x"397d5261",
1088 => x"5194f53f",
1089 => x"b00859b0",
1090 => x"08802e81",
1091 => x"a338b008",
1092 => x"f8056084",
1093 => x"0508fe06",
1094 => x"61055557",
1095 => x"76742e83",
1096 => x"e638fc18",
1097 => x"5675a426",
1098 => x"81aa387b",
1099 => x"b0085555",
1100 => x"93762780",
1101 => x"d8387470",
1102 => x"84055608",
1103 => x"b0087084",
1104 => x"05b00c0c",
1105 => x"b0087570",
1106 => x"84055708",
1107 => x"71708405",
1108 => x"530c549b",
1109 => x"7627b638",
1110 => x"74708405",
1111 => x"56087470",
1112 => x"8405560c",
1113 => x"74708405",
1114 => x"56087470",
1115 => x"8405560c",
1116 => x"a3762799",
1117 => x"38747084",
1118 => x"05560874",
1119 => x"70840556",
1120 => x"0c747084",
1121 => x"05560874",
1122 => x"70840556",
1123 => x"0c747084",
1124 => x"05560874",
1125 => x"70840556",
1126 => x"0c747084",
1127 => x"05560874",
1128 => x"70840556",
1129 => x"0c740874",
1130 => x"0c7b5261",
1131 => x"518bb83f",
1132 => x"6151a0ca",
1133 => x"3f785473",
1134 => x"b00c933d",
1135 => x"0d047d52",
1136 => x"615193b4",
1137 => x"3fb008b0",
1138 => x"0c933d0d",
1139 => x"04841608",
1140 => x"55fbd139",
1141 => x"75537b52",
1142 => x"b00851ef",
1143 => x"c83f7b52",
1144 => x"61518b83",
1145 => x"3fca398c",
1146 => x"16088817",
1147 => x"08718c12",
1148 => x"0c88120c",
1149 => x"558c1a08",
1150 => x"881b0871",
1151 => x"8c120c88",
1152 => x"120c5579",
1153 => x"795957fb",
1154 => x"f7397719",
1155 => x"901c5555",
1156 => x"737524fb",
1157 => x"a2387a17",
1158 => x"7080d984",
1159 => x"0b88050c",
1160 => x"757c3181",
1161 => x"0784120c",
1162 => x"5d841708",
1163 => x"81067b07",
1164 => x"84180c61",
1165 => x"519fc73f",
1166 => x"881754fc",
1167 => x"e5397419",
1168 => x"18901c55",
1169 => x"5d737d24",
1170 => x"fb95388c",
1171 => x"1a08881b",
1172 => x"08718c12",
1173 => x"0c88120c",
1174 => x"55881a61",
1175 => x"fc055759",
1176 => x"75a42681",
1177 => x"ae387b79",
1178 => x"55559376",
1179 => x"2780c938",
1180 => x"7b708405",
1181 => x"5d087c56",
1182 => x"790c7470",
1183 => x"84055608",
1184 => x"8c1b0c90",
1185 => x"1a549b76",
1186 => x"27ae3874",
1187 => x"70840556",
1188 => x"08740c74",
1189 => x"70840556",
1190 => x"08941b0c",
1191 => x"981a54a3",
1192 => x"76279538",
1193 => x"74708405",
1194 => x"5608740c",
1195 => x"74708405",
1196 => x"56089c1b",
1197 => x"0ca01a54",
1198 => x"74708405",
1199 => x"56087470",
1200 => x"8405560c",
1201 => x"74708405",
1202 => x"56087470",
1203 => x"8405560c",
1204 => x"7408740c",
1205 => x"7a1a7080",
1206 => x"d9840b88",
1207 => x"050c7d7c",
1208 => x"31810784",
1209 => x"120c5484",
1210 => x"1a088106",
1211 => x"7b07841b",
1212 => x"0c61519e",
1213 => x"893f7854",
1214 => x"fdbd3975",
1215 => x"537b5278",
1216 => x"51eda23f",
1217 => x"faf53984",
1218 => x"1708fc06",
1219 => x"18605858",
1220 => x"fae93975",
1221 => x"537b5278",
1222 => x"51ed8a3f",
1223 => x"7a1a7080",
1224 => x"d9840b88",
1225 => x"050c7d7c",
1226 => x"31810784",
1227 => x"120c5484",
1228 => x"1a088106",
1229 => x"7b07841b",
1230 => x"0cffb639",
1231 => x"fa3d0d78",
1232 => x"80d1c808",
1233 => x"5455b813",
1234 => x"08802e81",
1235 => x"b5388c15",
1236 => x"227083ff",
1237 => x"ff067083",
1238 => x"2a813270",
1239 => x"81065155",
1240 => x"55567280",
1241 => x"2e80dc38",
1242 => x"73842a81",
1243 => x"32810657",
1244 => x"ff537680",
1245 => x"f6387382",
1246 => x"2a708106",
1247 => x"51537280",
1248 => x"2eb938b0",
1249 => x"15085473",
1250 => x"802e9c38",
1251 => x"80c01553",
1252 => x"73732e8f",
1253 => x"38735280",
1254 => x"d1c80851",
1255 => x"87c93f8c",
1256 => x"15225676",
1257 => x"b0160c75",
1258 => x"db065372",
1259 => x"8c162380",
1260 => x"0b84160c",
1261 => x"90150875",
1262 => x"0c725675",
1263 => x"88075372",
1264 => x"8c162390",
1265 => x"1508802e",
1266 => x"80c0388c",
1267 => x"15227081",
1268 => x"06555373",
1269 => x"9d387281",
1270 => x"2a708106",
1271 => x"51537285",
1272 => x"38941508",
1273 => x"54738816",
1274 => x"0c805372",
1275 => x"b00c883d",
1276 => x"0d04800b",
1277 => x"88160c94",
1278 => x"15083098",
1279 => x"160c8053",
1280 => x"ea397251",
1281 => x"82fb3ffe",
1282 => x"c5397451",
1283 => x"8ce83f8c",
1284 => x"15227081",
1285 => x"06555373",
1286 => x"802effba",
1287 => x"38d439f8",
1288 => x"3d0d7a58",
1289 => x"77802e81",
1290 => x"993880d1",
1291 => x"c80854b8",
1292 => x"1408802e",
1293 => x"80ed388c",
1294 => x"18227090",
1295 => x"2b70902c",
1296 => x"70832a81",
1297 => x"3281065c",
1298 => x"51575478",
1299 => x"80cd3890",
1300 => x"18085776",
1301 => x"802e80c3",
1302 => x"38770877",
1303 => x"3177790c",
1304 => x"7683067a",
1305 => x"58555573",
1306 => x"85389418",
1307 => x"08567588",
1308 => x"190c8075",
1309 => x"25a53874",
1310 => x"5376529c",
1311 => x"180851a4",
1312 => x"18085473",
1313 => x"2d800bb0",
1314 => x"082580c9",
1315 => x"38b00817",
1316 => x"75b00831",
1317 => x"56577480",
1318 => x"24dd3880",
1319 => x"0bb00c8a",
1320 => x"3d0d0473",
1321 => x"5181da3f",
1322 => x"8c182270",
1323 => x"902b7090",
1324 => x"2c70832a",
1325 => x"81328106",
1326 => x"5c515754",
1327 => x"78dd38ff",
1328 => x"8e39a89f",
1329 => x"5280d1c8",
1330 => x"085189f1",
1331 => x"3fb008b0",
1332 => x"0c8a3d0d",
1333 => x"048c1822",
1334 => x"80c00754",
1335 => x"738c1923",
1336 => x"ff0bb00c",
1337 => x"8a3d0d04",
1338 => x"803d0d72",
1339 => x"5180710c",
1340 => x"800b8412",
1341 => x"0c800b88",
1342 => x"120c028e",
1343 => x"05228c12",
1344 => x"23029205",
1345 => x"228e1223",
1346 => x"800b9012",
1347 => x"0c800b94",
1348 => x"120c800b",
1349 => x"98120c70",
1350 => x"9c120c80",
1351 => x"c4b30ba0",
1352 => x"120c80c4",
1353 => x"ff0ba412",
1354 => x"0c80c5fb",
1355 => x"0ba8120c",
1356 => x"80c6cc0b",
1357 => x"ac120c82",
1358 => x"3d0d04fa",
1359 => x"3d0d7970",
1360 => x"80dc298c",
1361 => x"11547a53",
1362 => x"56578cac",
1363 => x"3fb008b0",
1364 => x"085556b0",
1365 => x"08802ea2",
1366 => x"38b0088c",
1367 => x"0554800b",
1368 => x"b0080c76",
1369 => x"b0088405",
1370 => x"0c73b008",
1371 => x"88050c74",
1372 => x"53805273",
1373 => x"5197f73f",
1374 => x"755473b0",
1375 => x"0c883d0d",
1376 => x"04fc3d0d",
1377 => x"76ad940b",
1378 => x"bc120c55",
1379 => x"810bb816",
1380 => x"0c800b84",
1381 => x"dc160c83",
1382 => x"0b84e016",
1383 => x"0c84e815",
1384 => x"84e4160c",
1385 => x"74548053",
1386 => x"84528415",
1387 => x"0851feb8",
1388 => x"3f745481",
1389 => x"53895288",
1390 => x"150851fe",
1391 => x"ab3f7454",
1392 => x"82538a52",
1393 => x"8c150851",
1394 => x"fe9e3f86",
1395 => x"3d0d04f9",
1396 => x"3d0d7980",
1397 => x"d1c80854",
1398 => x"57b81308",
1399 => x"802e80c8",
1400 => x"3884dc13",
1401 => x"56881608",
1402 => x"841708ff",
1403 => x"05555580",
1404 => x"74249f38",
1405 => x"8c152270",
1406 => x"902b7090",
1407 => x"2c515458",
1408 => x"72802e80",
1409 => x"ca3880dc",
1410 => x"15ff1555",
1411 => x"55738025",
1412 => x"e3387508",
1413 => x"5372802e",
1414 => x"9f387256",
1415 => x"88160884",
1416 => x"1708ff05",
1417 => x"5555c839",
1418 => x"7251fed5",
1419 => x"3f80d1c8",
1420 => x"0884dc05",
1421 => x"56ffae39",
1422 => x"84527651",
1423 => x"fdfd3fb0",
1424 => x"08760cb0",
1425 => x"08802e80",
1426 => x"c038b008",
1427 => x"56ce3981",
1428 => x"0b8c1623",
1429 => x"72750c72",
1430 => x"88160c72",
1431 => x"84160c72",
1432 => x"90160c72",
1433 => x"94160c72",
1434 => x"98160cff",
1435 => x"0b8e1623",
1436 => x"72b0160c",
1437 => x"72b4160c",
1438 => x"7280c416",
1439 => x"0c7280c8",
1440 => x"160c74b0",
1441 => x"0c893d0d",
1442 => x"048c770c",
1443 => x"800bb00c",
1444 => x"893d0d04",
1445 => x"ff3d0da8",
1446 => x"9f527351",
1447 => x"869f3f83",
1448 => x"3d0d0480",
1449 => x"3d0d80d1",
1450 => x"c80851e8",
1451 => x"3f823d0d",
1452 => x"04fb3d0d",
1453 => x"77705256",
1454 => x"96c33f80",
1455 => x"d9840b88",
1456 => x"05088411",
1457 => x"08fc0670",
1458 => x"7b319fef",
1459 => x"05e08006",
1460 => x"e0800556",
1461 => x"5653a080",
1462 => x"74249438",
1463 => x"80527551",
1464 => x"969d3f80",
1465 => x"d98c0815",
1466 => x"5372b008",
1467 => x"2e8f3875",
1468 => x"51968b3f",
1469 => x"805372b0",
1470 => x"0c873d0d",
1471 => x"04733052",
1472 => x"755195fb",
1473 => x"3fb008ff",
1474 => x"2ea83880",
1475 => x"d9840b88",
1476 => x"05087575",
1477 => x"31810784",
1478 => x"120c5380",
1479 => x"d8c80874",
1480 => x"3180d8c8",
1481 => x"0c755195",
1482 => x"d53f810b",
1483 => x"b00c873d",
1484 => x"0d048052",
1485 => x"755195c7",
1486 => x"3f80d984",
1487 => x"0b880508",
1488 => x"b0087131",
1489 => x"56538f75",
1490 => x"25ffa438",
1491 => x"b00880d8",
1492 => x"f8083180",
1493 => x"d8c80c74",
1494 => x"81078414",
1495 => x"0c755195",
1496 => x"9d3f8053",
1497 => x"ff9039f6",
1498 => x"3d0d7c7e",
1499 => x"545b7280",
1500 => x"2e828338",
1501 => x"7a519585",
1502 => x"3ff81384",
1503 => x"110870fe",
1504 => x"06701384",
1505 => x"1108fc06",
1506 => x"5d585954",
1507 => x"5880d98c",
1508 => x"08752e82",
1509 => x"de387884",
1510 => x"160c8073",
1511 => x"8106545a",
1512 => x"727a2e81",
1513 => x"d5387815",
1514 => x"84110881",
1515 => x"06515372",
1516 => x"a0387817",
1517 => x"577981e6",
1518 => x"38881508",
1519 => x"537280d9",
1520 => x"8c2e82f9",
1521 => x"388c1508",
1522 => x"708c150c",
1523 => x"7388120c",
1524 => x"56768107",
1525 => x"84190c76",
1526 => x"1877710c",
1527 => x"53798191",
1528 => x"3883ff77",
1529 => x"2781c838",
1530 => x"76892a77",
1531 => x"832a5653",
1532 => x"72802ebf",
1533 => x"3876862a",
1534 => x"b8055584",
1535 => x"7327b438",
1536 => x"80db1355",
1537 => x"947327ab",
1538 => x"38768c2a",
1539 => x"80ee0555",
1540 => x"80d47327",
1541 => x"9e38768f",
1542 => x"2a80f705",
1543 => x"5582d473",
1544 => x"27913876",
1545 => x"922a80fc",
1546 => x"05558ad4",
1547 => x"73278438",
1548 => x"80fe5574",
1549 => x"10101080",
1550 => x"d9840588",
1551 => x"11085556",
1552 => x"73762e82",
1553 => x"b3388414",
1554 => x"08fc0653",
1555 => x"7673278d",
1556 => x"38881408",
1557 => x"5473762e",
1558 => x"098106ea",
1559 => x"388c1408",
1560 => x"708c1a0c",
1561 => x"74881a0c",
1562 => x"7888120c",
1563 => x"56778c15",
1564 => x"0c7a5193",
1565 => x"893f8c3d",
1566 => x"0d047708",
1567 => x"78713159",
1568 => x"77058819",
1569 => x"08545772",
1570 => x"80d98c2e",
1571 => x"80e0388c",
1572 => x"1808708c",
1573 => x"150c7388",
1574 => x"120c56fe",
1575 => x"89398815",
1576 => x"088c1608",
1577 => x"708c130c",
1578 => x"5788170c",
1579 => x"fea33976",
1580 => x"832a7054",
1581 => x"55807524",
1582 => x"81983872",
1583 => x"822c8171",
1584 => x"2b80d988",
1585 => x"080780d9",
1586 => x"840b8405",
1587 => x"0c537410",
1588 => x"101080d9",
1589 => x"84058811",
1590 => x"08555675",
1591 => x"8c190c73",
1592 => x"88190c77",
1593 => x"88170c77",
1594 => x"8c150cff",
1595 => x"8439815a",
1596 => x"fdb43978",
1597 => x"17738106",
1598 => x"54577298",
1599 => x"38770878",
1600 => x"71315977",
1601 => x"058c1908",
1602 => x"881a0871",
1603 => x"8c120c88",
1604 => x"120c5757",
1605 => x"76810784",
1606 => x"190c7780",
1607 => x"d9840b88",
1608 => x"050c80d9",
1609 => x"80087726",
1610 => x"fec73880",
1611 => x"d8fc0852",
1612 => x"7a51fafd",
1613 => x"3f7a5191",
1614 => x"c53ffeba",
1615 => x"3981788c",
1616 => x"150c7888",
1617 => x"150c738c",
1618 => x"1a0c7388",
1619 => x"1a0c5afd",
1620 => x"80398315",
1621 => x"70822c81",
1622 => x"712b80d9",
1623 => x"88080780",
1624 => x"d9840b84",
1625 => x"050c5153",
1626 => x"74101010",
1627 => x"80d98405",
1628 => x"88110855",
1629 => x"56fee439",
1630 => x"74538075",
1631 => x"24a73872",
1632 => x"822c8171",
1633 => x"2b80d988",
1634 => x"080780d9",
1635 => x"840b8405",
1636 => x"0c53758c",
1637 => x"190c7388",
1638 => x"190c7788",
1639 => x"170c778c",
1640 => x"150cfdcd",
1641 => x"39831570",
1642 => x"822c8171",
1643 => x"2b80d988",
1644 => x"080780d9",
1645 => x"840b8405",
1646 => x"0c5153d6",
1647 => x"39f93d0d",
1648 => x"797b5853",
1649 => x"800b80d1",
1650 => x"c8085356",
1651 => x"72722e80",
1652 => x"c03884dc",
1653 => x"13557476",
1654 => x"2eb73888",
1655 => x"15088416",
1656 => x"08ff0554",
1657 => x"54807324",
1658 => x"9d388c14",
1659 => x"2270902b",
1660 => x"70902c51",
1661 => x"53587180",
1662 => x"d83880dc",
1663 => x"14ff1454",
1664 => x"54728025",
1665 => x"e5387408",
1666 => x"5574d038",
1667 => x"80d1c808",
1668 => x"5284dc12",
1669 => x"5574802e",
1670 => x"b1388815",
1671 => x"08841608",
1672 => x"ff055454",
1673 => x"8073249c",
1674 => x"388c1422",
1675 => x"70902b70",
1676 => x"902c5153",
1677 => x"5871ad38",
1678 => x"80dc14ff",
1679 => x"14545472",
1680 => x"8025e638",
1681 => x"74085574",
1682 => x"d13875b0",
1683 => x"0c893d0d",
1684 => x"04735176",
1685 => x"2d75b008",
1686 => x"0780dc15",
1687 => x"ff155555",
1688 => x"56ff9e39",
1689 => x"7351762d",
1690 => x"75b00807",
1691 => x"80dc15ff",
1692 => x"15555556",
1693 => x"ca39ea3d",
1694 => x"0d688c11",
1695 => x"2270812a",
1696 => x"81065758",
1697 => x"567480e4",
1698 => x"388e1622",
1699 => x"70902b70",
1700 => x"902c5155",
1701 => x"58807424",
1702 => x"b138983d",
1703 => x"c4055373",
1704 => x"5280d1c8",
1705 => x"085192ac",
1706 => x"3f800bb0",
1707 => x"08249738",
1708 => x"7983e080",
1709 => x"06547380",
1710 => x"c0802e81",
1711 => x"8f387382",
1712 => x"80802e81",
1713 => x"91388c16",
1714 => x"22577690",
1715 => x"80075473",
1716 => x"8c172388",
1717 => x"805280d1",
1718 => x"c8085181",
1719 => x"9b3fb008",
1720 => x"9d388c16",
1721 => x"22820754",
1722 => x"738c1723",
1723 => x"80c31670",
1724 => x"770c9017",
1725 => x"0c810b94",
1726 => x"170c983d",
1727 => x"0d0480d1",
1728 => x"c808ad94",
1729 => x"0bbc120c",
1730 => x"548c1622",
1731 => x"81800754",
1732 => x"738c1723",
1733 => x"b008760c",
1734 => x"b0089017",
1735 => x"0c88800b",
1736 => x"94170c74",
1737 => x"802ed338",
1738 => x"8e162270",
1739 => x"902b7090",
1740 => x"2c535558",
1741 => x"98ae3fb0",
1742 => x"08802eff",
1743 => x"bd388c16",
1744 => x"22810754",
1745 => x"738c1723",
1746 => x"983d0d04",
1747 => x"810b8c17",
1748 => x"225855fe",
1749 => x"f539a816",
1750 => x"0880c5fb",
1751 => x"2e098106",
1752 => x"fee4388c",
1753 => x"16228880",
1754 => x"0754738c",
1755 => x"17238880",
1756 => x"0b80cc17",
1757 => x"0cfedc39",
1758 => x"f33d0d7f",
1759 => x"618b1170",
1760 => x"f8065c55",
1761 => x"555e7296",
1762 => x"26833890",
1763 => x"59807924",
1764 => x"747a2607",
1765 => x"53805472",
1766 => x"742e0981",
1767 => x"0680cb38",
1768 => x"7d518cd9",
1769 => x"3f7883f7",
1770 => x"2680c638",
1771 => x"78832a70",
1772 => x"10101080",
1773 => x"d984058c",
1774 => x"11085959",
1775 => x"5a76782e",
1776 => x"83b03884",
1777 => x"1708fc06",
1778 => x"568c1708",
1779 => x"88180871",
1780 => x"8c120c88",
1781 => x"120c5875",
1782 => x"17841108",
1783 => x"81078412",
1784 => x"0c537d51",
1785 => x"8c983f88",
1786 => x"175473b0",
1787 => x"0c8f3d0d",
1788 => x"0478892a",
1789 => x"79832a5b",
1790 => x"5372802e",
1791 => x"bf387886",
1792 => x"2ab8055a",
1793 => x"847327b4",
1794 => x"3880db13",
1795 => x"5a947327",
1796 => x"ab38788c",
1797 => x"2a80ee05",
1798 => x"5a80d473",
1799 => x"279e3878",
1800 => x"8f2a80f7",
1801 => x"055a82d4",
1802 => x"73279138",
1803 => x"78922a80",
1804 => x"fc055a8a",
1805 => x"d4732784",
1806 => x"3880fe5a",
1807 => x"79101010",
1808 => x"80d98405",
1809 => x"8c110858",
1810 => x"5576752e",
1811 => x"a3388417",
1812 => x"08fc0670",
1813 => x"7a315556",
1814 => x"738f2488",
1815 => x"d5387380",
1816 => x"25fee638",
1817 => x"8c170857",
1818 => x"76752e09",
1819 => x"8106df38",
1820 => x"811a5a80",
1821 => x"d9940857",
1822 => x"7680d98c",
1823 => x"2e82c038",
1824 => x"841708fc",
1825 => x"06707a31",
1826 => x"5556738f",
1827 => x"2481f938",
1828 => x"80d98c0b",
1829 => x"80d9980c",
1830 => x"80d98c0b",
1831 => x"80d9940c",
1832 => x"738025fe",
1833 => x"b23883ff",
1834 => x"762783df",
1835 => x"3875892a",
1836 => x"76832a55",
1837 => x"5372802e",
1838 => x"bf387586",
1839 => x"2ab80554",
1840 => x"847327b4",
1841 => x"3880db13",
1842 => x"54947327",
1843 => x"ab38758c",
1844 => x"2a80ee05",
1845 => x"5480d473",
1846 => x"279e3875",
1847 => x"8f2a80f7",
1848 => x"055482d4",
1849 => x"73279138",
1850 => x"75922a80",
1851 => x"fc05548a",
1852 => x"d4732784",
1853 => x"3880fe54",
1854 => x"73101010",
1855 => x"80d98405",
1856 => x"88110856",
1857 => x"5874782e",
1858 => x"86cf3884",
1859 => x"1508fc06",
1860 => x"53757327",
1861 => x"8d388815",
1862 => x"08557478",
1863 => x"2e098106",
1864 => x"ea388c15",
1865 => x"0880d984",
1866 => x"0b840508",
1867 => x"718c1a0c",
1868 => x"76881a0c",
1869 => x"7888130c",
1870 => x"788c180c",
1871 => x"5d587953",
1872 => x"807a2483",
1873 => x"e6387282",
1874 => x"2c81712b",
1875 => x"5c537a7c",
1876 => x"26819838",
1877 => x"7b7b0653",
1878 => x"7282f138",
1879 => x"79fc0684",
1880 => x"055a7a10",
1881 => x"707d0654",
1882 => x"5b7282e0",
1883 => x"38841a5a",
1884 => x"f1398817",
1885 => x"8c110858",
1886 => x"5876782e",
1887 => x"098106fc",
1888 => x"c238821a",
1889 => x"5afdec39",
1890 => x"78177981",
1891 => x"0784190c",
1892 => x"7080d998",
1893 => x"0c7080d9",
1894 => x"940c80d9",
1895 => x"8c0b8c12",
1896 => x"0c8c1108",
1897 => x"88120c74",
1898 => x"81078412",
1899 => x"0c741175",
1900 => x"710c5153",
1901 => x"7d5188c6",
1902 => x"3f881754",
1903 => x"fcac3980",
1904 => x"d9840b84",
1905 => x"05087a54",
1906 => x"5c798025",
1907 => x"fef83882",
1908 => x"da397a09",
1909 => x"7c067080",
1910 => x"d9840b84",
1911 => x"050c5c7a",
1912 => x"105b7a7c",
1913 => x"2685387a",
1914 => x"85b83880",
1915 => x"d9840b88",
1916 => x"05087084",
1917 => x"1208fc06",
1918 => x"707c317c",
1919 => x"72268f72",
1920 => x"25075757",
1921 => x"5c5d5572",
1922 => x"802e80db",
1923 => x"38797a16",
1924 => x"80d8fc08",
1925 => x"1b90115a",
1926 => x"55575b80",
1927 => x"d8f808ff",
1928 => x"2e8838a0",
1929 => x"8f13e080",
1930 => x"06577652",
1931 => x"7d5187cf",
1932 => x"3fb00854",
1933 => x"b008ff2e",
1934 => x"9038b008",
1935 => x"76278299",
1936 => x"387480d9",
1937 => x"842e8291",
1938 => x"3880d984",
1939 => x"0b880508",
1940 => x"55841508",
1941 => x"fc06707a",
1942 => x"317a7226",
1943 => x"8f722507",
1944 => x"52555372",
1945 => x"83e63874",
1946 => x"79810784",
1947 => x"170c7916",
1948 => x"7080d984",
1949 => x"0b88050c",
1950 => x"75810784",
1951 => x"120c547e",
1952 => x"525786fa",
1953 => x"3f881754",
1954 => x"fae03975",
1955 => x"832a7054",
1956 => x"54807424",
1957 => x"819b3872",
1958 => x"822c8171",
1959 => x"2b80d988",
1960 => x"08077080",
1961 => x"d9840b84",
1962 => x"050c7510",
1963 => x"101080d9",
1964 => x"84058811",
1965 => x"08585a5d",
1966 => x"53778c18",
1967 => x"0c748818",
1968 => x"0c768819",
1969 => x"0c768c16",
1970 => x"0cfcf339",
1971 => x"797a1010",
1972 => x"1080d984",
1973 => x"05705759",
1974 => x"5d8c1508",
1975 => x"5776752e",
1976 => x"a3388417",
1977 => x"08fc0670",
1978 => x"7a315556",
1979 => x"738f2483",
1980 => x"ca387380",
1981 => x"25848138",
1982 => x"8c170857",
1983 => x"76752e09",
1984 => x"8106df38",
1985 => x"8815811b",
1986 => x"70830655",
1987 => x"5b5572c9",
1988 => x"387c8306",
1989 => x"5372802e",
1990 => x"fdb838ff",
1991 => x"1df81959",
1992 => x"5d881808",
1993 => x"782eea38",
1994 => x"fdb53983",
1995 => x"1a53fc96",
1996 => x"39831470",
1997 => x"822c8171",
1998 => x"2b80d988",
1999 => x"08077080",
2000 => x"d9840b84",
2001 => x"050c7610",
2002 => x"101080d9",
2003 => x"84058811",
2004 => x"08595b5e",
2005 => x"5153fee1",
2006 => x"3980d8c8",
2007 => x"081758b0",
2008 => x"08762e81",
2009 => x"8d3880d8",
2010 => x"f808ff2e",
2011 => x"83ec3873",
2012 => x"76311880",
2013 => x"d8c80c73",
2014 => x"87067057",
2015 => x"5372802e",
2016 => x"88388873",
2017 => x"31701555",
2018 => x"5676149f",
2019 => x"ff06a080",
2020 => x"71311770",
2021 => x"547f5357",
2022 => x"5384e43f",
2023 => x"b00853b0",
2024 => x"08ff2e81",
2025 => x"a03880d8",
2026 => x"c8081670",
2027 => x"80d8c80c",
2028 => x"747580d9",
2029 => x"840b8805",
2030 => x"0c747631",
2031 => x"18708107",
2032 => x"51555658",
2033 => x"7b80d984",
2034 => x"2e839c38",
2035 => x"798f2682",
2036 => x"cb38810b",
2037 => x"84150c84",
2038 => x"1508fc06",
2039 => x"707a317a",
2040 => x"72268f72",
2041 => x"25075255",
2042 => x"5372802e",
2043 => x"fcf93880",
2044 => x"db39b008",
2045 => x"9fff0653",
2046 => x"72feeb38",
2047 => x"7780d8c8",
2048 => x"0c80d984",
2049 => x"0b880508",
2050 => x"7b188107",
2051 => x"84120c55",
2052 => x"80d8f408",
2053 => x"78278638",
2054 => x"7780d8f4",
2055 => x"0c80d8f0",
2056 => x"087827fc",
2057 => x"ac387780",
2058 => x"d8f00c84",
2059 => x"1508fc06",
2060 => x"707a317a",
2061 => x"72268f72",
2062 => x"25075255",
2063 => x"5372802e",
2064 => x"fca53888",
2065 => x"39807454",
2066 => x"56fedb39",
2067 => x"7d5183ae",
2068 => x"3f800bb0",
2069 => x"0c8f3d0d",
2070 => x"04735380",
2071 => x"7424a938",
2072 => x"72822c81",
2073 => x"712b80d9",
2074 => x"88080770",
2075 => x"80d9840b",
2076 => x"84050c5d",
2077 => x"53778c18",
2078 => x"0c748818",
2079 => x"0c768819",
2080 => x"0c768c16",
2081 => x"0cf9b739",
2082 => x"83147082",
2083 => x"2c81712b",
2084 => x"80d98808",
2085 => x"077080d9",
2086 => x"840b8405",
2087 => x"0c5e5153",
2088 => x"d4397b7b",
2089 => x"065372fc",
2090 => x"a338841a",
2091 => x"7b105c5a",
2092 => x"f139ff1a",
2093 => x"8111515a",
2094 => x"f7b93978",
2095 => x"17798107",
2096 => x"84190c8c",
2097 => x"18088819",
2098 => x"08718c12",
2099 => x"0c88120c",
2100 => x"597080d9",
2101 => x"980c7080",
2102 => x"d9940c80",
2103 => x"d98c0b8c",
2104 => x"120c8c11",
2105 => x"0888120c",
2106 => x"74810784",
2107 => x"120c7411",
2108 => x"75710c51",
2109 => x"53f9bd39",
2110 => x"75178411",
2111 => x"08810784",
2112 => x"120c538c",
2113 => x"17088818",
2114 => x"08718c12",
2115 => x"0c88120c",
2116 => x"587d5181",
2117 => x"e93f8817",
2118 => x"54f5cf39",
2119 => x"7284150c",
2120 => x"f41af806",
2121 => x"70841e08",
2122 => x"81060784",
2123 => x"1e0c701d",
2124 => x"545b850b",
2125 => x"84140c85",
2126 => x"0b88140c",
2127 => x"8f7b27fd",
2128 => x"cf38881c",
2129 => x"527d51ec",
2130 => x"9e3f80d9",
2131 => x"840b8805",
2132 => x"0880d8c8",
2133 => x"085955fd",
2134 => x"b7397780",
2135 => x"d8c80c73",
2136 => x"80d8f80c",
2137 => x"fc913972",
2138 => x"84150cfd",
2139 => x"a339fc3d",
2140 => x"0d767971",
2141 => x"028c059f",
2142 => x"05335755",
2143 => x"53558372",
2144 => x"278a3874",
2145 => x"83065170",
2146 => x"802ea238",
2147 => x"ff125271",
2148 => x"ff2e9338",
2149 => x"73737081",
2150 => x"055534ff",
2151 => x"125271ff",
2152 => x"2e098106",
2153 => x"ef3874b0",
2154 => x"0c863d0d",
2155 => x"04747488",
2156 => x"2b750770",
2157 => x"71902b07",
2158 => x"5154518f",
2159 => x"7227a538",
2160 => x"72717084",
2161 => x"05530c72",
2162 => x"71708405",
2163 => x"530c7271",
2164 => x"70840553",
2165 => x"0c727170",
2166 => x"8405530c",
2167 => x"f0125271",
2168 => x"8f26dd38",
2169 => x"83722790",
2170 => x"38727170",
2171 => x"8405530c",
2172 => x"fc125271",
2173 => x"8326f238",
2174 => x"7053ff90",
2175 => x"390404fd",
2176 => x"3d0d800b",
2177 => x"80e1c00c",
2178 => x"765184ee",
2179 => x"3fb00853",
2180 => x"b008ff2e",
2181 => x"883872b0",
2182 => x"0c853d0d",
2183 => x"0480e1c0",
2184 => x"08547380",
2185 => x"2ef03875",
2186 => x"74710c52",
2187 => x"72b00c85",
2188 => x"3d0d04f9",
2189 => x"3d0d797c",
2190 => x"557b548e",
2191 => x"11227090",
2192 => x"2b70902c",
2193 => x"555780d1",
2194 => x"c8085358",
2195 => x"5683f33f",
2196 => x"b0085780",
2197 => x"0bb00824",
2198 => x"933880d0",
2199 => x"1608b008",
2200 => x"0580d017",
2201 => x"0c76b00c",
2202 => x"893d0d04",
2203 => x"8c162283",
2204 => x"dfff0655",
2205 => x"748c1723",
2206 => x"76b00c89",
2207 => x"3d0d04fa",
2208 => x"3d0d788c",
2209 => x"11227088",
2210 => x"2a708106",
2211 => x"51575856",
2212 => x"74a9388c",
2213 => x"162283df",
2214 => x"ff065574",
2215 => x"8c17237a",
2216 => x"5479538e",
2217 => x"16227090",
2218 => x"2b70902c",
2219 => x"545680d1",
2220 => x"c8085256",
2221 => x"81b23f88",
2222 => x"3d0d0482",
2223 => x"5480538e",
2224 => x"16227090",
2225 => x"2b70902c",
2226 => x"545680d1",
2227 => x"c8085257",
2228 => x"82b83f8c",
2229 => x"162283df",
2230 => x"ff065574",
2231 => x"8c17237a",
2232 => x"5479538e",
2233 => x"16227090",
2234 => x"2b70902c",
2235 => x"545680d1",
2236 => x"c8085256",
2237 => x"80f23f88",
2238 => x"3d0d04f9",
2239 => x"3d0d797c",
2240 => x"557b548e",
2241 => x"11227090",
2242 => x"2b70902c",
2243 => x"555780d1",
2244 => x"c8085358",
2245 => x"5681f33f",
2246 => x"b00857b0",
2247 => x"08ff2e99",
2248 => x"388c1622",
2249 => x"a0800755",
2250 => x"748c1723",
2251 => x"b00880d0",
2252 => x"170c76b0",
2253 => x"0c893d0d",
2254 => x"048c1622",
2255 => x"83dfff06",
2256 => x"55748c17",
2257 => x"2376b00c",
2258 => x"893d0d04",
2259 => x"fe3d0d74",
2260 => x"8e112270",
2261 => x"902b7090",
2262 => x"2c555151",
2263 => x"5380d1c8",
2264 => x"0851bd3f",
2265 => x"843d0d04",
2266 => x"fb3d0d80",
2267 => x"0b80e1c0",
2268 => x"0c7a5379",
2269 => x"52785182",
2270 => x"fb3fb008",
2271 => x"55b008ff",
2272 => x"2e883874",
2273 => x"b00c873d",
2274 => x"0d0480e1",
2275 => x"c0085675",
2276 => x"802ef038",
2277 => x"7776710c",
2278 => x"5474b00c",
2279 => x"873d0d04",
2280 => x"fd3d0d80",
2281 => x"0b80e1c0",
2282 => x"0c765184",
2283 => x"d03fb008",
2284 => x"53b008ff",
2285 => x"2e883872",
2286 => x"b00c853d",
2287 => x"0d0480e1",
2288 => x"c0085473",
2289 => x"802ef038",
2290 => x"7574710c",
2291 => x"5272b00c",
2292 => x"853d0d04",
2293 => x"fc3d0d80",
2294 => x"0b80e1c0",
2295 => x"0c785277",
2296 => x"5186b83f",
2297 => x"b00854b0",
2298 => x"08ff2e88",
2299 => x"3873b00c",
2300 => x"863d0d04",
2301 => x"80e1c008",
2302 => x"5574802e",
2303 => x"f0387675",
2304 => x"710c5373",
2305 => x"b00c863d",
2306 => x"0d04fb3d",
2307 => x"0d800b80",
2308 => x"e1c00c7a",
2309 => x"53795278",
2310 => x"5184943f",
2311 => x"b00855b0",
2312 => x"08ff2e88",
2313 => x"3874b00c",
2314 => x"873d0d04",
2315 => x"80e1c008",
2316 => x"5675802e",
2317 => x"f0387776",
2318 => x"710c5474",
2319 => x"b00c873d",
2320 => x"0d04fb3d",
2321 => x"0d800b80",
2322 => x"e1c00c7a",
2323 => x"53795278",
2324 => x"5182993f",
2325 => x"b00855b0",
2326 => x"08ff2e88",
2327 => x"3874b00c",
2328 => x"873d0d04",
2329 => x"80e1c008",
2330 => x"5675802e",
2331 => x"f0387776",
2332 => x"710c5474",
2333 => x"b00c873d",
2334 => x"0d04fe3d",
2335 => x"0d80e1b4",
2336 => x"0851708a",
2337 => x"3880e1c4",
2338 => x"7080e1b4",
2339 => x"0c517075",
2340 => x"125252ff",
2341 => x"537087fb",
2342 => x"80802688",
2343 => x"387080e1",
2344 => x"b40c7153",
2345 => x"72b00c84",
2346 => x"3d0d04fd",
2347 => x"3d0d800b",
2348 => x"80d1b808",
2349 => x"54547281",
2350 => x"2e9c3873",
2351 => x"80e1b80c",
2352 => x"c0a43fff",
2353 => x"beba3f80",
2354 => x"e18c5281",
2355 => x"51c2af3f",
2356 => x"b0085185",
2357 => x"c63f7280",
2358 => x"e1b80cc0",
2359 => x"893fffbe",
2360 => x"9f3f80e1",
2361 => x"8c528151",
2362 => x"c2943fb0",
2363 => x"085185ab",
2364 => x"3f00ff39",
2365 => x"f53d0d7e",
2366 => x"6080e1b8",
2367 => x"08705b58",
2368 => x"5b5b7580",
2369 => x"c538777a",
2370 => x"25a23877",
2371 => x"1b703370",
2372 => x"81ff0658",
2373 => x"5859758a",
2374 => x"2e993876",
2375 => x"81ff0651",
2376 => x"ffbfa23f",
2377 => x"81185879",
2378 => x"7824e038",
2379 => x"79b00c8d",
2380 => x"3d0d048d",
2381 => x"51ffbf8d",
2382 => x"3f783370",
2383 => x"81ff0652",
2384 => x"57ffbf81",
2385 => x"3f811858",
2386 => x"de397955",
2387 => x"7a547d53",
2388 => x"85528d3d",
2389 => x"fc0551ff",
2390 => x"bde83fb0",
2391 => x"085684b4",
2392 => x"3f7bb008",
2393 => x"0c75b00c",
2394 => x"8d3d0d04",
2395 => x"f63d0d7d",
2396 => x"7f80e1b8",
2397 => x"08705b58",
2398 => x"5a5a7580",
2399 => x"c4387779",
2400 => x"25b638ff",
2401 => x"be9a3fb0",
2402 => x"0881ff06",
2403 => x"708d3270",
2404 => x"30709f2a",
2405 => x"51515757",
2406 => x"768a2e80",
2407 => x"c6387580",
2408 => x"2e80c038",
2409 => x"771a5676",
2410 => x"76347651",
2411 => x"ffbe963f",
2412 => x"81185878",
2413 => x"7824cc38",
2414 => x"775675b0",
2415 => x"0c8c3d0d",
2416 => x"04785579",
2417 => x"547c5384",
2418 => x"528c3dfc",
2419 => x"0551ffbc",
2420 => x"f13fb008",
2421 => x"5683bd3f",
2422 => x"7ab0080c",
2423 => x"75b00c8c",
2424 => x"3d0d0477",
2425 => x"1a568a76",
2426 => x"34811858",
2427 => x"8d51ffbd",
2428 => x"d43f8a51",
2429 => x"ffbdce3f",
2430 => x"7756ffbe",
2431 => x"39fb3d0d",
2432 => x"80e1b808",
2433 => x"70565473",
2434 => x"883874b0",
2435 => x"0c873d0d",
2436 => x"04775383",
2437 => x"52873dfc",
2438 => x"0551ffbc",
2439 => x"a53fb008",
2440 => x"5482f13f",
2441 => x"75b0080c",
2442 => x"73b00c87",
2443 => x"3d0d04fa",
2444 => x"3d0d80e1",
2445 => x"b808802e",
2446 => x"a3387a55",
2447 => x"79547853",
2448 => x"8652883d",
2449 => x"fc0551ff",
2450 => x"bbf83fb0",
2451 => x"085682c4",
2452 => x"3f76b008",
2453 => x"0c75b00c",
2454 => x"883d0d04",
2455 => x"82b63f9d",
2456 => x"0bb0080c",
2457 => x"ff0bb00c",
2458 => x"883d0d04",
2459 => x"fb3d0d77",
2460 => x"79565680",
2461 => x"70545473",
2462 => x"75259f38",
2463 => x"74101010",
2464 => x"f8055272",
2465 => x"16703370",
2466 => x"742b7607",
2467 => x"8116f816",
2468 => x"56565651",
2469 => x"51747324",
2470 => x"ea3873b0",
2471 => x"0c873d0d",
2472 => x"04fc3d0d",
2473 => x"76785555",
2474 => x"bc538052",
2475 => x"7351f5be",
2476 => x"3f845274",
2477 => x"51ffb53f",
2478 => x"b0087423",
2479 => x"84528415",
2480 => x"51ffa93f",
2481 => x"b0088215",
2482 => x"23845288",
2483 => x"1551ff9c",
2484 => x"3fb00884",
2485 => x"150c8452",
2486 => x"8c1551ff",
2487 => x"8f3fb008",
2488 => x"88152384",
2489 => x"52901551",
2490 => x"ff823fb0",
2491 => x"088a1523",
2492 => x"84529415",
2493 => x"51fef53f",
2494 => x"b0088c15",
2495 => x"23845298",
2496 => x"1551fee8",
2497 => x"3fb0088e",
2498 => x"15238852",
2499 => x"9c1551fe",
2500 => x"db3fb008",
2501 => x"90150c86",
2502 => x"3d0d04e9",
2503 => x"3d0d6a80",
2504 => x"e1b80857",
2505 => x"57759338",
2506 => x"80c0800b",
2507 => x"84180c75",
2508 => x"ac180c75",
2509 => x"b00c993d",
2510 => x"0d04893d",
2511 => x"70556a54",
2512 => x"558a5299",
2513 => x"3dffbc05",
2514 => x"51ffb9f6",
2515 => x"3fb00877",
2516 => x"53755256",
2517 => x"fecb3fbc",
2518 => x"3f77b008",
2519 => x"0c75b00c",
2520 => x"993d0d04",
2521 => x"fc3d0d81",
2522 => x"5480e1b8",
2523 => x"08883873",
2524 => x"b00c863d",
2525 => x"0d047653",
2526 => x"97b95286",
2527 => x"3dfc0551",
2528 => x"ffb9bf3f",
2529 => x"b008548c",
2530 => x"3f74b008",
2531 => x"0c73b00c",
2532 => x"863d0d04",
2533 => x"80d1c808",
2534 => x"b00c04f7",
2535 => x"3d0d7b80",
2536 => x"d1c80882",
2537 => x"c811085a",
2538 => x"545a7780",
2539 => x"2e80da38",
2540 => x"81881884",
2541 => x"1908ff05",
2542 => x"81712b59",
2543 => x"55598074",
2544 => x"2480ea38",
2545 => x"807424b5",
2546 => x"3873822b",
2547 => x"78118805",
2548 => x"56568180",
2549 => x"19087706",
2550 => x"5372802e",
2551 => x"b6387816",
2552 => x"70085353",
2553 => x"79517408",
2554 => x"53722dff",
2555 => x"14fc17fc",
2556 => x"1779812c",
2557 => x"5a575754",
2558 => x"738025d6",
2559 => x"38770858",
2560 => x"77ffad38",
2561 => x"80d1c808",
2562 => x"53bc1308",
2563 => x"a5387951",
2564 => x"f9df3f74",
2565 => x"0853722d",
2566 => x"ff14fc17",
2567 => x"fc177981",
2568 => x"2c5a5757",
2569 => x"54738025",
2570 => x"ffa838d1",
2571 => x"398057ff",
2572 => x"93397251",
2573 => x"bc130853",
2574 => x"722d7951",
2575 => x"f9b33fff",
2576 => x"3d0d80e1",
2577 => x"940bfc05",
2578 => x"70085252",
2579 => x"70ff2e91",
2580 => x"38702dfc",
2581 => x"12700852",
2582 => x"5270ff2e",
2583 => x"098106f1",
2584 => x"38833d0d",
2585 => x"0404ffb9",
2586 => x"e83f0400",
2587 => x"00ffffff",
2588 => x"ff00ffff",
2589 => x"ffff00ff",
2590 => x"ffffff00",
2591 => x"00000040",
2592 => x"30313233",
2593 => x"34353637",
2594 => x"38396162",
2595 => x"63646566",
2596 => x"00000000",
2597 => x"633a0000",
2598 => x"733a0000",
2599 => x"623a0000",
2600 => x"0a000000",
2601 => x"43000000",
2602 => x"64756d6d",
2603 => x"792e6578",
2604 => x"65000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"0000309c",
2609 => x"00002880",
2610 => x"000028cc",
2611 => x"00000000",
2612 => x"00002b34",
2613 => x"00002b90",
2614 => x"00002bec",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"000028a4",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000001",
2654 => x"330eabcd",
2655 => x"1234e66d",
2656 => x"deec0005",
2657 => x"000b0000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000000",
2827 => x"00000000",
2828 => x"00000000",
2829 => x"00000000",
2830 => x"00000000",
2831 => x"00000000",
2832 => x"00000000",
2833 => x"00000000",
2834 => x"00000000",
2835 => x"00000000",
2836 => x"00000000",
2837 => x"00000000",
2838 => x"00000000",
2839 => x"00000000",
2840 => x"00000000",
2841 => x"00000000",
2842 => x"00000000",
2843 => x"00000000",
2844 => x"00000000",
2845 => x"00000000",
2846 => x"ffffffff",
2847 => x"00000000",
2848 => x"00020000",
2849 => x"00000000",
2850 => x"00000000",
2851 => x"00002c84",
2852 => x"00002c84",
2853 => x"00002c8c",
2854 => x"00002c8c",
2855 => x"00002c94",
2856 => x"00002c94",
2857 => x"00002c9c",
2858 => x"00002c9c",
2859 => x"00002ca4",
2860 => x"00002ca4",
2861 => x"00002cac",
2862 => x"00002cac",
2863 => x"00002cb4",
2864 => x"00002cb4",
2865 => x"00002cbc",
2866 => x"00002cbc",
2867 => x"00002cc4",
2868 => x"00002cc4",
2869 => x"00002ccc",
2870 => x"00002ccc",
2871 => x"00002cd4",
2872 => x"00002cd4",
2873 => x"00002cdc",
2874 => x"00002cdc",
2875 => x"00002ce4",
2876 => x"00002ce4",
2877 => x"00002cec",
2878 => x"00002cec",
2879 => x"00002cf4",
2880 => x"00002cf4",
2881 => x"00002cfc",
2882 => x"00002cfc",
2883 => x"00002d04",
2884 => x"00002d04",
2885 => x"00002d0c",
2886 => x"00002d0c",
2887 => x"00002d14",
2888 => x"00002d14",
2889 => x"00002d1c",
2890 => x"00002d1c",
2891 => x"00002d24",
2892 => x"00002d24",
2893 => x"00002d2c",
2894 => x"00002d2c",
2895 => x"00002d34",
2896 => x"00002d34",
2897 => x"00002d3c",
2898 => x"00002d3c",
2899 => x"00002d44",
2900 => x"00002d44",
2901 => x"00002d4c",
2902 => x"00002d4c",
2903 => x"00002d54",
2904 => x"00002d54",
2905 => x"00002d5c",
2906 => x"00002d5c",
2907 => x"00002d64",
2908 => x"00002d64",
2909 => x"00002d6c",
2910 => x"00002d6c",
2911 => x"00002d74",
2912 => x"00002d74",
2913 => x"00002d7c",
2914 => x"00002d7c",
2915 => x"00002d84",
2916 => x"00002d84",
2917 => x"00002d8c",
2918 => x"00002d8c",
2919 => x"00002d94",
2920 => x"00002d94",
2921 => x"00002d9c",
2922 => x"00002d9c",
2923 => x"00002da4",
2924 => x"00002da4",
2925 => x"00002dac",
2926 => x"00002dac",
2927 => x"00002db4",
2928 => x"00002db4",
2929 => x"00002dbc",
2930 => x"00002dbc",
2931 => x"00002dc4",
2932 => x"00002dc4",
2933 => x"00002dcc",
2934 => x"00002dcc",
2935 => x"00002dd4",
2936 => x"00002dd4",
2937 => x"00002ddc",
2938 => x"00002ddc",
2939 => x"00002de4",
2940 => x"00002de4",
2941 => x"00002dec",
2942 => x"00002dec",
2943 => x"00002df4",
2944 => x"00002df4",
2945 => x"00002dfc",
2946 => x"00002dfc",
2947 => x"00002e04",
2948 => x"00002e04",
2949 => x"00002e0c",
2950 => x"00002e0c",
2951 => x"00002e14",
2952 => x"00002e14",
2953 => x"00002e1c",
2954 => x"00002e1c",
2955 => x"00002e24",
2956 => x"00002e24",
2957 => x"00002e2c",
2958 => x"00002e2c",
2959 => x"00002e34",
2960 => x"00002e34",
2961 => x"00002e3c",
2962 => x"00002e3c",
2963 => x"00002e44",
2964 => x"00002e44",
2965 => x"00002e4c",
2966 => x"00002e4c",
2967 => x"00002e54",
2968 => x"00002e54",
2969 => x"00002e5c",
2970 => x"00002e5c",
2971 => x"00002e64",
2972 => x"00002e64",
2973 => x"00002e6c",
2974 => x"00002e6c",
2975 => x"00002e74",
2976 => x"00002e74",
2977 => x"00002e7c",
2978 => x"00002e7c",
2979 => x"00002e84",
2980 => x"00002e84",
2981 => x"00002e8c",
2982 => x"00002e8c",
2983 => x"00002e94",
2984 => x"00002e94",
2985 => x"00002e9c",
2986 => x"00002e9c",
2987 => x"00002ea4",
2988 => x"00002ea4",
2989 => x"00002eac",
2990 => x"00002eac",
2991 => x"00002eb4",
2992 => x"00002eb4",
2993 => x"00002ebc",
2994 => x"00002ebc",
2995 => x"00002ec4",
2996 => x"00002ec4",
2997 => x"00002ecc",
2998 => x"00002ecc",
2999 => x"00002ed4",
3000 => x"00002ed4",
3001 => x"00002edc",
3002 => x"00002edc",
3003 => x"00002ee4",
3004 => x"00002ee4",
3005 => x"00002eec",
3006 => x"00002eec",
3007 => x"00002ef4",
3008 => x"00002ef4",
3009 => x"00002efc",
3010 => x"00002efc",
3011 => x"00002f04",
3012 => x"00002f04",
3013 => x"00002f0c",
3014 => x"00002f0c",
3015 => x"00002f14",
3016 => x"00002f14",
3017 => x"00002f1c",
3018 => x"00002f1c",
3019 => x"00002f24",
3020 => x"00002f24",
3021 => x"00002f2c",
3022 => x"00002f2c",
3023 => x"00002f34",
3024 => x"00002f34",
3025 => x"00002f3c",
3026 => x"00002f3c",
3027 => x"00002f44",
3028 => x"00002f44",
3029 => x"00002f4c",
3030 => x"00002f4c",
3031 => x"00002f54",
3032 => x"00002f54",
3033 => x"00002f5c",
3034 => x"00002f5c",
3035 => x"00002f64",
3036 => x"00002f64",
3037 => x"00002f6c",
3038 => x"00002f6c",
3039 => x"00002f74",
3040 => x"00002f74",
3041 => x"00002f7c",
3042 => x"00002f7c",
3043 => x"00002f84",
3044 => x"00002f84",
3045 => x"00002f8c",
3046 => x"00002f8c",
3047 => x"00002f94",
3048 => x"00002f94",
3049 => x"00002f9c",
3050 => x"00002f9c",
3051 => x"00002fa4",
3052 => x"00002fa4",
3053 => x"00002fac",
3054 => x"00002fac",
3055 => x"00002fb4",
3056 => x"00002fb4",
3057 => x"00002fbc",
3058 => x"00002fbc",
3059 => x"00002fc4",
3060 => x"00002fc4",
3061 => x"00002fcc",
3062 => x"00002fcc",
3063 => x"00002fd4",
3064 => x"00002fd4",
3065 => x"00002fdc",
3066 => x"00002fdc",
3067 => x"00002fe4",
3068 => x"00002fe4",
3069 => x"00002fec",
3070 => x"00002fec",
3071 => x"00002ff4",
3072 => x"00002ff4",
3073 => x"00002ffc",
3074 => x"00002ffc",
3075 => x"00003004",
3076 => x"00003004",
3077 => x"0000300c",
3078 => x"0000300c",
3079 => x"00003014",
3080 => x"00003014",
3081 => x"0000301c",
3082 => x"0000301c",
3083 => x"00003024",
3084 => x"00003024",
3085 => x"0000302c",
3086 => x"0000302c",
3087 => x"00003034",
3088 => x"00003034",
3089 => x"0000303c",
3090 => x"0000303c",
3091 => x"00003044",
3092 => x"00003044",
3093 => x"0000304c",
3094 => x"0000304c",
3095 => x"00003054",
3096 => x"00003054",
3097 => x"0000305c",
3098 => x"0000305c",
3099 => x"00003064",
3100 => x"00003064",
3101 => x"0000306c",
3102 => x"0000306c",
3103 => x"00003074",
3104 => x"00003074",
3105 => x"0000307c",
3106 => x"0000307c",
3107 => x"000028a8",
3108 => x"ffffffff",
3109 => x"00000000",
3110 => x"ffffffff",
3111 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

