------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cdf00c",
3 => x"3a0b0b80",
4 => x"c5f50400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80cd",
162 => x"a8738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cdec0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c4f63f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8da32d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8bf12d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80ddd8",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80dd",
307 => x"d8085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480cd",
314 => x"ec08802e",
315 => x"a43880cd",
316 => x"f008822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80ddd80c",
320 => x"82a0800b",
321 => x"80dddc0c",
322 => x"8290800b",
323 => x"80dde00c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80ddd8",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"dddc0cf8",
330 => x"80808480",
331 => x"0b80dde0",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80dd",
335 => x"d80c80c0",
336 => x"a880940b",
337 => x"80dddc0c",
338 => x"80cdb80b",
339 => x"80dde00c",
340 => x"04ff3d0d",
341 => x"80dde433",
342 => x"5170a738",
343 => x"80cdf808",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"cdf80c70",
348 => x"2d80cdf8",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80dd",
352 => x"e434833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80ddd408",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"ddd4510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404803d",
366 => x"0d80ddf0",
367 => x"08811180",
368 => x"ddf00c51",
369 => x"823d0d04",
370 => x"fe3d0d80",
371 => x"ddf00853",
372 => x"80ddf008",
373 => x"5272722e",
374 => x"8f3880cd",
375 => x"bc5185e8",
376 => x"3f80ddf0",
377 => x"0853e939",
378 => x"80cdcc51",
379 => x"85da3fe0",
380 => x"39bc0802",
381 => x"bc0cf93d",
382 => x"0d800bbc",
383 => x"08fc050c",
384 => x"bc088805",
385 => x"088025ab",
386 => x"38bc0888",
387 => x"050830bc",
388 => x"0888050c",
389 => x"800bbc08",
390 => x"f4050cbc",
391 => x"08fc0508",
392 => x"8838810b",
393 => x"bc08f405",
394 => x"0cbc08f4",
395 => x"0508bc08",
396 => x"fc050cbc",
397 => x"088c0508",
398 => x"8025ab38",
399 => x"bc088c05",
400 => x"0830bc08",
401 => x"8c050c80",
402 => x"0bbc08f0",
403 => x"050cbc08",
404 => x"fc050888",
405 => x"38810bbc",
406 => x"08f0050c",
407 => x"bc08f005",
408 => x"08bc08fc",
409 => x"050c8053",
410 => x"bc088c05",
411 => x"0852bc08",
412 => x"88050851",
413 => x"81a73fb0",
414 => x"0870bc08",
415 => x"f8050c54",
416 => x"bc08fc05",
417 => x"08802e8c",
418 => x"38bc08f8",
419 => x"050830bc",
420 => x"08f8050c",
421 => x"bc08f805",
422 => x"0870b00c",
423 => x"54893d0d",
424 => x"bc0c04bc",
425 => x"0802bc0c",
426 => x"fb3d0d80",
427 => x"0bbc08fc",
428 => x"050cbc08",
429 => x"88050880",
430 => x"259338bc",
431 => x"08880508",
432 => x"30bc0888",
433 => x"050c810b",
434 => x"bc08fc05",
435 => x"0cbc088c",
436 => x"05088025",
437 => x"8c38bc08",
438 => x"8c050830",
439 => x"bc088c05",
440 => x"0c8153bc",
441 => x"088c0508",
442 => x"52bc0888",
443 => x"050851ad",
444 => x"3fb00870",
445 => x"bc08f805",
446 => x"0c54bc08",
447 => x"fc050880",
448 => x"2e8c38bc",
449 => x"08f80508",
450 => x"30bc08f8",
451 => x"050cbc08",
452 => x"f8050870",
453 => x"b00c5487",
454 => x"3d0dbc0c",
455 => x"04bc0802",
456 => x"bc0cfd3d",
457 => x"0d810bbc",
458 => x"08fc050c",
459 => x"800bbc08",
460 => x"f8050cbc",
461 => x"088c0508",
462 => x"bc088805",
463 => x"0827ac38",
464 => x"bc08fc05",
465 => x"08802ea3",
466 => x"38800bbc",
467 => x"088c0508",
468 => x"249938bc",
469 => x"088c0508",
470 => x"10bc088c",
471 => x"050cbc08",
472 => x"fc050810",
473 => x"bc08fc05",
474 => x"0cc939bc",
475 => x"08fc0508",
476 => x"802e80c9",
477 => x"38bc088c",
478 => x"0508bc08",
479 => x"88050826",
480 => x"a138bc08",
481 => x"880508bc",
482 => x"088c0508",
483 => x"31bc0888",
484 => x"050cbc08",
485 => x"f80508bc",
486 => x"08fc0508",
487 => x"07bc08f8",
488 => x"050cbc08",
489 => x"fc050881",
490 => x"2abc08fc",
491 => x"050cbc08",
492 => x"8c050881",
493 => x"2abc088c",
494 => x"050cffaf",
495 => x"39bc0890",
496 => x"0508802e",
497 => x"8f38bc08",
498 => x"88050870",
499 => x"bc08f405",
500 => x"0c518d39",
501 => x"bc08f805",
502 => x"0870bc08",
503 => x"f4050c51",
504 => x"bc08f405",
505 => x"08b00c85",
506 => x"3d0dbc0c",
507 => x"04fc3d0d",
508 => x"7670797b",
509 => x"55555555",
510 => x"8f72278c",
511 => x"38727507",
512 => x"83065170",
513 => x"802ea738",
514 => x"ff125271",
515 => x"ff2e9838",
516 => x"72708105",
517 => x"54337470",
518 => x"81055634",
519 => x"ff125271",
520 => x"ff2e0981",
521 => x"06ea3874",
522 => x"b00c863d",
523 => x"0d047451",
524 => x"72708405",
525 => x"54087170",
526 => x"8405530c",
527 => x"72708405",
528 => x"54087170",
529 => x"8405530c",
530 => x"72708405",
531 => x"54087170",
532 => x"8405530c",
533 => x"72708405",
534 => x"54087170",
535 => x"8405530c",
536 => x"f0125271",
537 => x"8f26c938",
538 => x"83722795",
539 => x"38727084",
540 => x"05540871",
541 => x"70840553",
542 => x"0cfc1252",
543 => x"718326ed",
544 => x"387054ff",
545 => x"8339f73d",
546 => x"0d7c7052",
547 => x"5380ca3f",
548 => x"7254b008",
549 => x"550b0b80",
550 => x"cdd85681",
551 => x"57b00881",
552 => x"055a8b3d",
553 => x"e4115953",
554 => x"8259f413",
555 => x"527b8811",
556 => x"08525381",
557 => x"833fb008",
558 => x"3070b008",
559 => x"079f2c8a",
560 => x"07b00c53",
561 => x"8b3d0d04",
562 => x"ff3d0d73",
563 => x"5280cdfc",
564 => x"0851ffb2",
565 => x"3f833d0d",
566 => x"04fd3d0d",
567 => x"75707183",
568 => x"06535552",
569 => x"70b83871",
570 => x"70087009",
571 => x"f7fbfdff",
572 => x"120670f8",
573 => x"84828180",
574 => x"06515152",
575 => x"53709d38",
576 => x"84137008",
577 => x"7009f7fb",
578 => x"fdff1206",
579 => x"70f88482",
580 => x"81800651",
581 => x"51525370",
582 => x"802ee538",
583 => x"72527133",
584 => x"5170802e",
585 => x"8a388112",
586 => x"70335252",
587 => x"70f83871",
588 => x"7431b00c",
589 => x"853d0d04",
590 => x"f23d0d60",
591 => x"62881108",
592 => x"7057575f",
593 => x"5a74802e",
594 => x"818f388c",
595 => x"1a227083",
596 => x"2a813270",
597 => x"81065155",
598 => x"58738638",
599 => x"901a0891",
600 => x"38795190",
601 => x"a13fff54",
602 => x"b00880ed",
603 => x"388c1a22",
604 => x"587d0857",
605 => x"807883ff",
606 => x"ff067081",
607 => x"2a708106",
608 => x"51565755",
609 => x"73752e80",
610 => x"d7387490",
611 => x"38760884",
612 => x"18088819",
613 => x"59565974",
614 => x"802ef238",
615 => x"74548880",
616 => x"75278438",
617 => x"88805473",
618 => x"5378529c",
619 => x"1a0851a4",
620 => x"1a085473",
621 => x"2d800bb0",
622 => x"082582e6",
623 => x"38b00819",
624 => x"75b00831",
625 => x"7f880508",
626 => x"b0083170",
627 => x"6188050c",
628 => x"56565973",
629 => x"ffb43880",
630 => x"5473b00c",
631 => x"903d0d04",
632 => x"75813270",
633 => x"81067641",
634 => x"51547380",
635 => x"2e81c138",
636 => x"74903876",
637 => x"08841808",
638 => x"88195956",
639 => x"5974802e",
640 => x"f238881a",
641 => x"087883ff",
642 => x"ff067089",
643 => x"2a708106",
644 => x"51565956",
645 => x"73802e82",
646 => x"fa387575",
647 => x"278d3877",
648 => x"872a7081",
649 => x"06515473",
650 => x"82b53874",
651 => x"76278338",
652 => x"74567553",
653 => x"78527908",
654 => x"5185823f",
655 => x"881a0876",
656 => x"31881b0c",
657 => x"7908167a",
658 => x"0c745675",
659 => x"19757731",
660 => x"7f880508",
661 => x"78317061",
662 => x"88050c56",
663 => x"56597380",
664 => x"2efef438",
665 => x"8c1a2258",
666 => x"ff863977",
667 => x"78547953",
668 => x"7b525684",
669 => x"c83f881a",
670 => x"08783188",
671 => x"1b0c7908",
672 => x"187a0c7c",
673 => x"76315d7c",
674 => x"8e387951",
675 => x"8fdb3fb0",
676 => x"08818f38",
677 => x"b0085f75",
678 => x"19757731",
679 => x"7f880508",
680 => x"78317061",
681 => x"88050c56",
682 => x"56597380",
683 => x"2efea838",
684 => x"74818338",
685 => x"76088418",
686 => x"08881959",
687 => x"56597480",
688 => x"2ef23874",
689 => x"538a5278",
690 => x"5182d33f",
691 => x"b0087931",
692 => x"81055db0",
693 => x"08843881",
694 => x"155d815f",
695 => x"7c58747d",
696 => x"27833874",
697 => x"58941a08",
698 => x"881b0811",
699 => x"575c807a",
700 => x"085c5490",
701 => x"1a087b27",
702 => x"83388154",
703 => x"75782584",
704 => x"3873ba38",
705 => x"7b7824fe",
706 => x"e2387b53",
707 => x"78529c1a",
708 => x"0851a41a",
709 => x"0854732d",
710 => x"b00856b0",
711 => x"088024fe",
712 => x"e2388c1a",
713 => x"2280c007",
714 => x"54738c1b",
715 => x"23ff5473",
716 => x"b00c903d",
717 => x"0d047eff",
718 => x"a338ff87",
719 => x"39755378",
720 => x"527a5182",
721 => x"f83f7908",
722 => x"167a0c79",
723 => x"518e9a3f",
724 => x"b008cf38",
725 => x"7c76315d",
726 => x"7cfebc38",
727 => x"feac3990",
728 => x"1a087a08",
729 => x"71317611",
730 => x"70565a57",
731 => x"5280cdfc",
732 => x"0851848c",
733 => x"3fb00880",
734 => x"2effa738",
735 => x"b008901b",
736 => x"0cb00816",
737 => x"7a0c7794",
738 => x"1b0c7488",
739 => x"1b0c7456",
740 => x"fd993979",
741 => x"0858901a",
742 => x"08782783",
743 => x"38815475",
744 => x"75278438",
745 => x"73b33894",
746 => x"1a085675",
747 => x"752680d3",
748 => x"38755378",
749 => x"529c1a08",
750 => x"51a41a08",
751 => x"54732db0",
752 => x"0856b008",
753 => x"8024fd83",
754 => x"388c1a22",
755 => x"80c00754",
756 => x"738c1b23",
757 => x"ff54fed7",
758 => x"39755378",
759 => x"52775181",
760 => x"dc3f7908",
761 => x"167a0c79",
762 => x"518cfe3f",
763 => x"b008802e",
764 => x"fcd9388c",
765 => x"1a2280c0",
766 => x"0754738c",
767 => x"1b23ff54",
768 => x"fead3974",
769 => x"75547953",
770 => x"78525681",
771 => x"b03f881a",
772 => x"08753188",
773 => x"1b0c7908",
774 => x"157a0cfc",
775 => x"ae39fa3d",
776 => x"0d7a7902",
777 => x"8805a705",
778 => x"33565253",
779 => x"8373278a",
780 => x"38708306",
781 => x"5271802e",
782 => x"a838ff13",
783 => x"5372ff2e",
784 => x"97387033",
785 => x"5273722e",
786 => x"91388111",
787 => x"ff145451",
788 => x"72ff2e09",
789 => x"8106eb38",
790 => x"805170b0",
791 => x"0c883d0d",
792 => x"04707257",
793 => x"55835175",
794 => x"82802914",
795 => x"ff125256",
796 => x"708025f3",
797 => x"38837327",
798 => x"bf387408",
799 => x"76327009",
800 => x"f7fbfdff",
801 => x"120670f8",
802 => x"84828180",
803 => x"06515151",
804 => x"70802e99",
805 => x"38745180",
806 => x"52703357",
807 => x"73772eff",
808 => x"b9388111",
809 => x"81135351",
810 => x"837227ed",
811 => x"38fc1384",
812 => x"16565372",
813 => x"8326c338",
814 => x"7451fefe",
815 => x"39fa3d0d",
816 => x"787a7c72",
817 => x"72725757",
818 => x"57595656",
819 => x"747627b2",
820 => x"38761551",
821 => x"757127aa",
822 => x"38707717",
823 => x"ff145455",
824 => x"5371ff2e",
825 => x"9638ff14",
826 => x"ff145454",
827 => x"72337434",
828 => x"ff125271",
829 => x"ff2e0981",
830 => x"06ec3875",
831 => x"b00c883d",
832 => x"0d04768f",
833 => x"269738ff",
834 => x"125271ff",
835 => x"2eed3872",
836 => x"70810554",
837 => x"33747081",
838 => x"055634eb",
839 => x"39747607",
840 => x"83065170",
841 => x"e2387575",
842 => x"54517270",
843 => x"84055408",
844 => x"71708405",
845 => x"530c7270",
846 => x"84055408",
847 => x"71708405",
848 => x"530c7270",
849 => x"84055408",
850 => x"71708405",
851 => x"530c7270",
852 => x"84055408",
853 => x"71708405",
854 => x"530cf012",
855 => x"52718f26",
856 => x"c9388372",
857 => x"27953872",
858 => x"70840554",
859 => x"08717084",
860 => x"05530cfc",
861 => x"12527183",
862 => x"26ed3870",
863 => x"54ff8839",
864 => x"ef3d0d63",
865 => x"6567405d",
866 => x"427b802e",
867 => x"84fa3861",
868 => x"51a5b43f",
869 => x"f81c7084",
870 => x"120870fc",
871 => x"0670628b",
872 => x"0570f806",
873 => x"4159455b",
874 => x"5c415796",
875 => x"742782c3",
876 => x"38807b24",
877 => x"7e7c2607",
878 => x"59805478",
879 => x"742e0981",
880 => x"0682a938",
881 => x"777b2581",
882 => x"fc387717",
883 => x"80d5b80b",
884 => x"8805085e",
885 => x"567c762e",
886 => x"84bd3884",
887 => x"160870fe",
888 => x"06178411",
889 => x"08810651",
890 => x"55557382",
891 => x"8b3874fc",
892 => x"06597c76",
893 => x"2e84dd38",
894 => x"77195f7e",
895 => x"7b2581fd",
896 => x"38798106",
897 => x"547382bf",
898 => x"38767708",
899 => x"31841108",
900 => x"fc06565a",
901 => x"75802e91",
902 => x"387c762e",
903 => x"84ea3874",
904 => x"19185978",
905 => x"7b258489",
906 => x"3879802e",
907 => x"82993877",
908 => x"15567a76",
909 => x"24829038",
910 => x"8c1a0888",
911 => x"1b08718c",
912 => x"120c8812",
913 => x"0c557976",
914 => x"59578817",
915 => x"61fc0557",
916 => x"5975a426",
917 => x"85ef387b",
918 => x"79555593",
919 => x"762780c9",
920 => x"387b7084",
921 => x"055d087c",
922 => x"56790c74",
923 => x"70840556",
924 => x"088c180c",
925 => x"9017549b",
926 => x"7627ae38",
927 => x"74708405",
928 => x"5608740c",
929 => x"74708405",
930 => x"56089418",
931 => x"0c981754",
932 => x"a3762795",
933 => x"38747084",
934 => x"05560874",
935 => x"0c747084",
936 => x"0556089c",
937 => x"180ca017",
938 => x"54747084",
939 => x"05560874",
940 => x"70840556",
941 => x"0c747084",
942 => x"05560874",
943 => x"70840556",
944 => x"0c740874",
945 => x"0c777b31",
946 => x"56758f26",
947 => x"80c93884",
948 => x"17088106",
949 => x"78078418",
950 => x"0c771784",
951 => x"11088107",
952 => x"84120c54",
953 => x"6151a2e0",
954 => x"3f881754",
955 => x"73b00c93",
956 => x"3d0d0490",
957 => x"5bfdba39",
958 => x"7856fe85",
959 => x"398c1608",
960 => x"88170871",
961 => x"8c120c88",
962 => x"120c557e",
963 => x"707c3157",
964 => x"588f7627",
965 => x"ffb9387a",
966 => x"17841808",
967 => x"81067c07",
968 => x"84190c76",
969 => x"81078412",
970 => x"0c761184",
971 => x"11088107",
972 => x"84120c55",
973 => x"88055261",
974 => x"518cf63f",
975 => x"6151a288",
976 => x"3f881754",
977 => x"ffa6397d",
978 => x"52615194",
979 => x"f53fb008",
980 => x"59b00880",
981 => x"2e81a338",
982 => x"b008f805",
983 => x"60840508",
984 => x"fe066105",
985 => x"55577674",
986 => x"2e83e638",
987 => x"fc185675",
988 => x"a42681aa",
989 => x"387bb008",
990 => x"55559376",
991 => x"2780d838",
992 => x"74708405",
993 => x"5608b008",
994 => x"708405b0",
995 => x"0c0cb008",
996 => x"75708405",
997 => x"57087170",
998 => x"8405530c",
999 => x"549b7627",
1000 => x"b6387470",
1001 => x"84055608",
1002 => x"74708405",
1003 => x"560c7470",
1004 => x"84055608",
1005 => x"74708405",
1006 => x"560ca376",
1007 => x"27993874",
1008 => x"70840556",
1009 => x"08747084",
1010 => x"05560c74",
1011 => x"70840556",
1012 => x"08747084",
1013 => x"05560c74",
1014 => x"70840556",
1015 => x"08747084",
1016 => x"05560c74",
1017 => x"70840556",
1018 => x"08747084",
1019 => x"05560c74",
1020 => x"08740c7b",
1021 => x"5261518b",
1022 => x"b83f6151",
1023 => x"a0ca3f78",
1024 => x"5473b00c",
1025 => x"933d0d04",
1026 => x"7d526151",
1027 => x"93b43fb0",
1028 => x"08b00c93",
1029 => x"3d0d0484",
1030 => x"160855fb",
1031 => x"d1397553",
1032 => x"7b52b008",
1033 => x"51efc63f",
1034 => x"7b526151",
1035 => x"8b833fca",
1036 => x"398c1608",
1037 => x"88170871",
1038 => x"8c120c88",
1039 => x"120c558c",
1040 => x"1a08881b",
1041 => x"08718c12",
1042 => x"0c88120c",
1043 => x"55797959",
1044 => x"57fbf739",
1045 => x"7719901c",
1046 => x"55557375",
1047 => x"24fba238",
1048 => x"7a177080",
1049 => x"d5b80b88",
1050 => x"050c757c",
1051 => x"31810784",
1052 => x"120c5d84",
1053 => x"17088106",
1054 => x"7b078418",
1055 => x"0c61519f",
1056 => x"c73f8817",
1057 => x"54fce539",
1058 => x"74191890",
1059 => x"1c555d73",
1060 => x"7d24fb95",
1061 => x"388c1a08",
1062 => x"881b0871",
1063 => x"8c120c88",
1064 => x"120c5588",
1065 => x"1a61fc05",
1066 => x"575975a4",
1067 => x"2681ae38",
1068 => x"7b795555",
1069 => x"93762780",
1070 => x"c9387b70",
1071 => x"84055d08",
1072 => x"7c56790c",
1073 => x"74708405",
1074 => x"56088c1b",
1075 => x"0c901a54",
1076 => x"9b7627ae",
1077 => x"38747084",
1078 => x"05560874",
1079 => x"0c747084",
1080 => x"05560894",
1081 => x"1b0c981a",
1082 => x"54a37627",
1083 => x"95387470",
1084 => x"84055608",
1085 => x"740c7470",
1086 => x"84055608",
1087 => x"9c1b0ca0",
1088 => x"1a547470",
1089 => x"84055608",
1090 => x"74708405",
1091 => x"560c7470",
1092 => x"84055608",
1093 => x"74708405",
1094 => x"560c7408",
1095 => x"740c7a1a",
1096 => x"7080d5b8",
1097 => x"0b88050c",
1098 => x"7d7c3181",
1099 => x"0784120c",
1100 => x"54841a08",
1101 => x"81067b07",
1102 => x"841b0c61",
1103 => x"519e893f",
1104 => x"7854fdbd",
1105 => x"3975537b",
1106 => x"527851ed",
1107 => x"a03ffaf5",
1108 => x"39841708",
1109 => x"fc061860",
1110 => x"5858fae9",
1111 => x"3975537b",
1112 => x"527851ed",
1113 => x"883f7a1a",
1114 => x"7080d5b8",
1115 => x"0b88050c",
1116 => x"7d7c3181",
1117 => x"0784120c",
1118 => x"54841a08",
1119 => x"81067b07",
1120 => x"841b0cff",
1121 => x"b639fa3d",
1122 => x"0d7880cd",
1123 => x"fc085455",
1124 => x"b8130880",
1125 => x"2e81b538",
1126 => x"8c152270",
1127 => x"83ffff06",
1128 => x"70832a81",
1129 => x"32708106",
1130 => x"51555556",
1131 => x"72802e80",
1132 => x"dc387384",
1133 => x"2a813281",
1134 => x"0657ff53",
1135 => x"7680f638",
1136 => x"73822a70",
1137 => x"81065153",
1138 => x"72802eb9",
1139 => x"38b01508",
1140 => x"5473802e",
1141 => x"9c3880c0",
1142 => x"15537373",
1143 => x"2e8f3873",
1144 => x"5280cdfc",
1145 => x"085187c9",
1146 => x"3f8c1522",
1147 => x"5676b016",
1148 => x"0c75db06",
1149 => x"53728c16",
1150 => x"23800b84",
1151 => x"160c9015",
1152 => x"08750c72",
1153 => x"56758807",
1154 => x"53728c16",
1155 => x"23901508",
1156 => x"802e80c0",
1157 => x"388c1522",
1158 => x"70810655",
1159 => x"53739d38",
1160 => x"72812a70",
1161 => x"81065153",
1162 => x"72853894",
1163 => x"15085473",
1164 => x"88160c80",
1165 => x"5372b00c",
1166 => x"883d0d04",
1167 => x"800b8816",
1168 => x"0c941508",
1169 => x"3098160c",
1170 => x"8053ea39",
1171 => x"725182fb",
1172 => x"3ffec539",
1173 => x"74518ce8",
1174 => x"3f8c1522",
1175 => x"70810655",
1176 => x"5373802e",
1177 => x"ffba38d4",
1178 => x"39f83d0d",
1179 => x"7a587780",
1180 => x"2e819938",
1181 => x"80cdfc08",
1182 => x"54b81408",
1183 => x"802e80ed",
1184 => x"388c1822",
1185 => x"70902b70",
1186 => x"902c7083",
1187 => x"2a813281",
1188 => x"065c5157",
1189 => x"547880cd",
1190 => x"38901808",
1191 => x"5776802e",
1192 => x"80c33877",
1193 => x"08773177",
1194 => x"790c7683",
1195 => x"067a5855",
1196 => x"55738538",
1197 => x"94180856",
1198 => x"7588190c",
1199 => x"807525a5",
1200 => x"38745376",
1201 => x"529c1808",
1202 => x"51a41808",
1203 => x"54732d80",
1204 => x"0bb00825",
1205 => x"80c938b0",
1206 => x"081775b0",
1207 => x"08315657",
1208 => x"748024dd",
1209 => x"38800bb0",
1210 => x"0c8a3d0d",
1211 => x"04735181",
1212 => x"da3f8c18",
1213 => x"2270902b",
1214 => x"70902c70",
1215 => x"832a8132",
1216 => x"81065c51",
1217 => x"575478dd",
1218 => x"38ff8e39",
1219 => x"a4e95280",
1220 => x"cdfc0851",
1221 => x"89f13fb0",
1222 => x"08b00c8a",
1223 => x"3d0d048c",
1224 => x"182280c0",
1225 => x"0754738c",
1226 => x"1923ff0b",
1227 => x"b00c8a3d",
1228 => x"0d04803d",
1229 => x"0d725180",
1230 => x"710c800b",
1231 => x"84120c80",
1232 => x"0b88120c",
1233 => x"028e0522",
1234 => x"8c122302",
1235 => x"9205228e",
1236 => x"1223800b",
1237 => x"90120c80",
1238 => x"0b94120c",
1239 => x"800b9812",
1240 => x"0c709c12",
1241 => x"0c80c0fd",
1242 => x"0ba0120c",
1243 => x"80c1c90b",
1244 => x"a4120c80",
1245 => x"c2c50ba8",
1246 => x"120c80c3",
1247 => x"960bac12",
1248 => x"0c823d0d",
1249 => x"04fa3d0d",
1250 => x"797080dc",
1251 => x"298c1154",
1252 => x"7a535657",
1253 => x"8cac3fb0",
1254 => x"08b00855",
1255 => x"56b00880",
1256 => x"2ea238b0",
1257 => x"088c0554",
1258 => x"800bb008",
1259 => x"0c76b008",
1260 => x"84050c73",
1261 => x"b0088805",
1262 => x"0c745380",
1263 => x"52735197",
1264 => x"f73f7554",
1265 => x"73b00c88",
1266 => x"3d0d04fc",
1267 => x"3d0d76a9",
1268 => x"de0bbc12",
1269 => x"0c55810b",
1270 => x"b8160c80",
1271 => x"0b84dc16",
1272 => x"0c830b84",
1273 => x"e0160c84",
1274 => x"e81584e4",
1275 => x"160c7454",
1276 => x"80538452",
1277 => x"84150851",
1278 => x"feb83f74",
1279 => x"54815389",
1280 => x"52881508",
1281 => x"51feab3f",
1282 => x"74548253",
1283 => x"8a528c15",
1284 => x"0851fe9e",
1285 => x"3f863d0d",
1286 => x"04f93d0d",
1287 => x"7980cdfc",
1288 => x"085457b8",
1289 => x"1308802e",
1290 => x"80c83884",
1291 => x"dc135688",
1292 => x"16088417",
1293 => x"08ff0555",
1294 => x"55807424",
1295 => x"9f388c15",
1296 => x"2270902b",
1297 => x"70902c51",
1298 => x"54587280",
1299 => x"2e80ca38",
1300 => x"80dc15ff",
1301 => x"15555573",
1302 => x"8025e338",
1303 => x"75085372",
1304 => x"802e9f38",
1305 => x"72568816",
1306 => x"08841708",
1307 => x"ff055555",
1308 => x"c8397251",
1309 => x"fed53f80",
1310 => x"cdfc0884",
1311 => x"dc0556ff",
1312 => x"ae398452",
1313 => x"7651fdfd",
1314 => x"3fb00876",
1315 => x"0cb00880",
1316 => x"2e80c038",
1317 => x"b00856ce",
1318 => x"39810b8c",
1319 => x"16237275",
1320 => x"0c728816",
1321 => x"0c728416",
1322 => x"0c729016",
1323 => x"0c729416",
1324 => x"0c729816",
1325 => x"0cff0b8e",
1326 => x"162372b0",
1327 => x"160c72b4",
1328 => x"160c7280",
1329 => x"c4160c72",
1330 => x"80c8160c",
1331 => x"74b00c89",
1332 => x"3d0d048c",
1333 => x"770c800b",
1334 => x"b00c893d",
1335 => x"0d04ff3d",
1336 => x"0da4e952",
1337 => x"7351869f",
1338 => x"3f833d0d",
1339 => x"04803d0d",
1340 => x"80cdfc08",
1341 => x"51e83f82",
1342 => x"3d0d04fb",
1343 => x"3d0d7770",
1344 => x"525696c3",
1345 => x"3f80d5b8",
1346 => x"0b880508",
1347 => x"841108fc",
1348 => x"06707b31",
1349 => x"9fef05e0",
1350 => x"8006e080",
1351 => x"05565653",
1352 => x"a0807424",
1353 => x"94388052",
1354 => x"7551969d",
1355 => x"3f80d5c0",
1356 => x"08155372",
1357 => x"b0082e8f",
1358 => x"38755196",
1359 => x"8b3f8053",
1360 => x"72b00c87",
1361 => x"3d0d0473",
1362 => x"30527551",
1363 => x"95fb3fb0",
1364 => x"08ff2ea8",
1365 => x"3880d5b8",
1366 => x"0b880508",
1367 => x"75753181",
1368 => x"0784120c",
1369 => x"5380d4fc",
1370 => x"08743180",
1371 => x"d4fc0c75",
1372 => x"5195d53f",
1373 => x"810bb00c",
1374 => x"873d0d04",
1375 => x"80527551",
1376 => x"95c73f80",
1377 => x"d5b80b88",
1378 => x"0508b008",
1379 => x"71315653",
1380 => x"8f7525ff",
1381 => x"a438b008",
1382 => x"80d5ac08",
1383 => x"3180d4fc",
1384 => x"0c748107",
1385 => x"84140c75",
1386 => x"51959d3f",
1387 => x"8053ff90",
1388 => x"39f63d0d",
1389 => x"7c7e545b",
1390 => x"72802e82",
1391 => x"83387a51",
1392 => x"95853ff8",
1393 => x"13841108",
1394 => x"70fe0670",
1395 => x"13841108",
1396 => x"fc065d58",
1397 => x"59545880",
1398 => x"d5c00875",
1399 => x"2e82de38",
1400 => x"7884160c",
1401 => x"80738106",
1402 => x"545a727a",
1403 => x"2e81d538",
1404 => x"78158411",
1405 => x"08810651",
1406 => x"5372a038",
1407 => x"78175779",
1408 => x"81e63888",
1409 => x"15085372",
1410 => x"80d5c02e",
1411 => x"82f9388c",
1412 => x"1508708c",
1413 => x"150c7388",
1414 => x"120c5676",
1415 => x"81078419",
1416 => x"0c761877",
1417 => x"710c5379",
1418 => x"81913883",
1419 => x"ff772781",
1420 => x"c8387689",
1421 => x"2a77832a",
1422 => x"56537280",
1423 => x"2ebf3876",
1424 => x"862ab805",
1425 => x"55847327",
1426 => x"b43880db",
1427 => x"13559473",
1428 => x"27ab3876",
1429 => x"8c2a80ee",
1430 => x"055580d4",
1431 => x"73279e38",
1432 => x"768f2a80",
1433 => x"f7055582",
1434 => x"d4732791",
1435 => x"3876922a",
1436 => x"80fc0555",
1437 => x"8ad47327",
1438 => x"843880fe",
1439 => x"55741010",
1440 => x"1080d5b8",
1441 => x"05881108",
1442 => x"55567376",
1443 => x"2e82b338",
1444 => x"841408fc",
1445 => x"06537673",
1446 => x"278d3888",
1447 => x"14085473",
1448 => x"762e0981",
1449 => x"06ea388c",
1450 => x"1408708c",
1451 => x"1a0c7488",
1452 => x"1a0c7888",
1453 => x"120c5677",
1454 => x"8c150c7a",
1455 => x"5193893f",
1456 => x"8c3d0d04",
1457 => x"77087871",
1458 => x"31597705",
1459 => x"88190854",
1460 => x"577280d5",
1461 => x"c02e80e0",
1462 => x"388c1808",
1463 => x"708c150c",
1464 => x"7388120c",
1465 => x"56fe8939",
1466 => x"8815088c",
1467 => x"1608708c",
1468 => x"130c5788",
1469 => x"170cfea3",
1470 => x"3976832a",
1471 => x"70545580",
1472 => x"75248198",
1473 => x"3872822c",
1474 => x"81712b80",
1475 => x"d5bc0807",
1476 => x"80d5b80b",
1477 => x"84050c53",
1478 => x"74101010",
1479 => x"80d5b805",
1480 => x"88110855",
1481 => x"56758c19",
1482 => x"0c738819",
1483 => x"0c778817",
1484 => x"0c778c15",
1485 => x"0cff8439",
1486 => x"815afdb4",
1487 => x"39781773",
1488 => x"81065457",
1489 => x"72983877",
1490 => x"08787131",
1491 => x"5977058c",
1492 => x"1908881a",
1493 => x"08718c12",
1494 => x"0c88120c",
1495 => x"57577681",
1496 => x"0784190c",
1497 => x"7780d5b8",
1498 => x"0b88050c",
1499 => x"80d5b408",
1500 => x"7726fec7",
1501 => x"3880d5b0",
1502 => x"08527a51",
1503 => x"fafd3f7a",
1504 => x"5191c53f",
1505 => x"feba3981",
1506 => x"788c150c",
1507 => x"7888150c",
1508 => x"738c1a0c",
1509 => x"73881a0c",
1510 => x"5afd8039",
1511 => x"83157082",
1512 => x"2c81712b",
1513 => x"80d5bc08",
1514 => x"0780d5b8",
1515 => x"0b84050c",
1516 => x"51537410",
1517 => x"101080d5",
1518 => x"b8058811",
1519 => x"085556fe",
1520 => x"e4397453",
1521 => x"807524a7",
1522 => x"3872822c",
1523 => x"81712b80",
1524 => x"d5bc0807",
1525 => x"80d5b80b",
1526 => x"84050c53",
1527 => x"758c190c",
1528 => x"7388190c",
1529 => x"7788170c",
1530 => x"778c150c",
1531 => x"fdcd3983",
1532 => x"1570822c",
1533 => x"81712b80",
1534 => x"d5bc0807",
1535 => x"80d5b80b",
1536 => x"84050c51",
1537 => x"53d639f9",
1538 => x"3d0d797b",
1539 => x"5853800b",
1540 => x"80cdfc08",
1541 => x"53567272",
1542 => x"2e80c038",
1543 => x"84dc1355",
1544 => x"74762eb7",
1545 => x"38881508",
1546 => x"841608ff",
1547 => x"05545480",
1548 => x"73249d38",
1549 => x"8c142270",
1550 => x"902b7090",
1551 => x"2c515358",
1552 => x"7180d838",
1553 => x"80dc14ff",
1554 => x"14545472",
1555 => x"8025e538",
1556 => x"74085574",
1557 => x"d03880cd",
1558 => x"fc085284",
1559 => x"dc125574",
1560 => x"802eb138",
1561 => x"88150884",
1562 => x"1608ff05",
1563 => x"54548073",
1564 => x"249c388c",
1565 => x"14227090",
1566 => x"2b70902c",
1567 => x"51535871",
1568 => x"ad3880dc",
1569 => x"14ff1454",
1570 => x"54728025",
1571 => x"e6387408",
1572 => x"5574d138",
1573 => x"75b00c89",
1574 => x"3d0d0473",
1575 => x"51762d75",
1576 => x"b0080780",
1577 => x"dc15ff15",
1578 => x"555556ff",
1579 => x"9e397351",
1580 => x"762d75b0",
1581 => x"080780dc",
1582 => x"15ff1555",
1583 => x"5556ca39",
1584 => x"ea3d0d68",
1585 => x"8c112270",
1586 => x"812a8106",
1587 => x"57585674",
1588 => x"80e4388e",
1589 => x"16227090",
1590 => x"2b70902c",
1591 => x"51555880",
1592 => x"7424b138",
1593 => x"983dc405",
1594 => x"53735280",
1595 => x"cdfc0851",
1596 => x"92ac3f80",
1597 => x"0bb00824",
1598 => x"97387983",
1599 => x"e0800654",
1600 => x"7380c080",
1601 => x"2e818f38",
1602 => x"73828080",
1603 => x"2e819138",
1604 => x"8c162257",
1605 => x"76908007",
1606 => x"54738c17",
1607 => x"23888052",
1608 => x"80cdfc08",
1609 => x"51819b3f",
1610 => x"b0089d38",
1611 => x"8c162282",
1612 => x"0754738c",
1613 => x"172380c3",
1614 => x"1670770c",
1615 => x"90170c81",
1616 => x"0b94170c",
1617 => x"983d0d04",
1618 => x"80cdfc08",
1619 => x"a9de0bbc",
1620 => x"120c548c",
1621 => x"16228180",
1622 => x"0754738c",
1623 => x"1723b008",
1624 => x"760cb008",
1625 => x"90170c88",
1626 => x"800b9417",
1627 => x"0c74802e",
1628 => x"d3388e16",
1629 => x"2270902b",
1630 => x"70902c53",
1631 => x"555898a1",
1632 => x"3fb00880",
1633 => x"2effbd38",
1634 => x"8c162281",
1635 => x"0754738c",
1636 => x"1723983d",
1637 => x"0d04810b",
1638 => x"8c172258",
1639 => x"55fef539",
1640 => x"a8160880",
1641 => x"c2c52e09",
1642 => x"8106fee4",
1643 => x"388c1622",
1644 => x"88800754",
1645 => x"738c1723",
1646 => x"88800b80",
1647 => x"cc170cfe",
1648 => x"dc39f33d",
1649 => x"0d7f618b",
1650 => x"1170f806",
1651 => x"5c55555e",
1652 => x"72962683",
1653 => x"38905980",
1654 => x"7924747a",
1655 => x"26075380",
1656 => x"5472742e",
1657 => x"09810680",
1658 => x"cb387d51",
1659 => x"8cd93f78",
1660 => x"83f72680",
1661 => x"c6387883",
1662 => x"2a701010",
1663 => x"1080d5b8",
1664 => x"058c1108",
1665 => x"59595a76",
1666 => x"782e83b0",
1667 => x"38841708",
1668 => x"fc06568c",
1669 => x"17088818",
1670 => x"08718c12",
1671 => x"0c88120c",
1672 => x"58751784",
1673 => x"11088107",
1674 => x"84120c53",
1675 => x"7d518c98",
1676 => x"3f881754",
1677 => x"73b00c8f",
1678 => x"3d0d0478",
1679 => x"892a7983",
1680 => x"2a5b5372",
1681 => x"802ebf38",
1682 => x"78862ab8",
1683 => x"055a8473",
1684 => x"27b43880",
1685 => x"db135a94",
1686 => x"7327ab38",
1687 => x"788c2a80",
1688 => x"ee055a80",
1689 => x"d473279e",
1690 => x"38788f2a",
1691 => x"80f7055a",
1692 => x"82d47327",
1693 => x"91387892",
1694 => x"2a80fc05",
1695 => x"5a8ad473",
1696 => x"27843880",
1697 => x"fe5a7910",
1698 => x"101080d5",
1699 => x"b8058c11",
1700 => x"08585576",
1701 => x"752ea338",
1702 => x"841708fc",
1703 => x"06707a31",
1704 => x"5556738f",
1705 => x"2488d538",
1706 => x"738025fe",
1707 => x"e6388c17",
1708 => x"08577675",
1709 => x"2e098106",
1710 => x"df38811a",
1711 => x"5a80d5c8",
1712 => x"08577680",
1713 => x"d5c02e82",
1714 => x"c0388417",
1715 => x"08fc0670",
1716 => x"7a315556",
1717 => x"738f2481",
1718 => x"f93880d5",
1719 => x"c00b80d5",
1720 => x"cc0c80d5",
1721 => x"c00b80d5",
1722 => x"c80c7380",
1723 => x"25feb238",
1724 => x"83ff7627",
1725 => x"83df3875",
1726 => x"892a7683",
1727 => x"2a555372",
1728 => x"802ebf38",
1729 => x"75862ab8",
1730 => x"05548473",
1731 => x"27b43880",
1732 => x"db135494",
1733 => x"7327ab38",
1734 => x"758c2a80",
1735 => x"ee055480",
1736 => x"d473279e",
1737 => x"38758f2a",
1738 => x"80f70554",
1739 => x"82d47327",
1740 => x"91387592",
1741 => x"2a80fc05",
1742 => x"548ad473",
1743 => x"27843880",
1744 => x"fe547310",
1745 => x"101080d5",
1746 => x"b8058811",
1747 => x"08565874",
1748 => x"782e86cf",
1749 => x"38841508",
1750 => x"fc065375",
1751 => x"73278d38",
1752 => x"88150855",
1753 => x"74782e09",
1754 => x"8106ea38",
1755 => x"8c150880",
1756 => x"d5b80b84",
1757 => x"0508718c",
1758 => x"1a0c7688",
1759 => x"1a0c7888",
1760 => x"130c788c",
1761 => x"180c5d58",
1762 => x"7953807a",
1763 => x"2483e638",
1764 => x"72822c81",
1765 => x"712b5c53",
1766 => x"7a7c2681",
1767 => x"98387b7b",
1768 => x"06537282",
1769 => x"f13879fc",
1770 => x"0684055a",
1771 => x"7a10707d",
1772 => x"06545b72",
1773 => x"82e03884",
1774 => x"1a5af139",
1775 => x"88178c11",
1776 => x"08585876",
1777 => x"782e0981",
1778 => x"06fcc238",
1779 => x"821a5afd",
1780 => x"ec397817",
1781 => x"79810784",
1782 => x"190c7080",
1783 => x"d5cc0c70",
1784 => x"80d5c80c",
1785 => x"80d5c00b",
1786 => x"8c120c8c",
1787 => x"11088812",
1788 => x"0c748107",
1789 => x"84120c74",
1790 => x"1175710c",
1791 => x"51537d51",
1792 => x"88c63f88",
1793 => x"1754fcac",
1794 => x"3980d5b8",
1795 => x"0b840508",
1796 => x"7a545c79",
1797 => x"8025fef8",
1798 => x"3882da39",
1799 => x"7a097c06",
1800 => x"7080d5b8",
1801 => x"0b84050c",
1802 => x"5c7a105b",
1803 => x"7a7c2685",
1804 => x"387a85b8",
1805 => x"3880d5b8",
1806 => x"0b880508",
1807 => x"70841208",
1808 => x"fc06707c",
1809 => x"317c7226",
1810 => x"8f722507",
1811 => x"57575c5d",
1812 => x"5572802e",
1813 => x"80db3879",
1814 => x"7a1680d5",
1815 => x"b0081b90",
1816 => x"115a5557",
1817 => x"5b80d5ac",
1818 => x"08ff2e88",
1819 => x"38a08f13",
1820 => x"e0800657",
1821 => x"76527d51",
1822 => x"87cf3fb0",
1823 => x"0854b008",
1824 => x"ff2e9038",
1825 => x"b0087627",
1826 => x"82993874",
1827 => x"80d5b82e",
1828 => x"82913880",
1829 => x"d5b80b88",
1830 => x"05085584",
1831 => x"1508fc06",
1832 => x"707a317a",
1833 => x"72268f72",
1834 => x"25075255",
1835 => x"537283e6",
1836 => x"38747981",
1837 => x"0784170c",
1838 => x"79167080",
1839 => x"d5b80b88",
1840 => x"050c7581",
1841 => x"0784120c",
1842 => x"547e5257",
1843 => x"86fa3f88",
1844 => x"1754fae0",
1845 => x"3975832a",
1846 => x"70545480",
1847 => x"7424819b",
1848 => x"3872822c",
1849 => x"81712b80",
1850 => x"d5bc0807",
1851 => x"7080d5b8",
1852 => x"0b84050c",
1853 => x"75101010",
1854 => x"80d5b805",
1855 => x"88110858",
1856 => x"5a5d5377",
1857 => x"8c180c74",
1858 => x"88180c76",
1859 => x"88190c76",
1860 => x"8c160cfc",
1861 => x"f339797a",
1862 => x"10101080",
1863 => x"d5b80570",
1864 => x"57595d8c",
1865 => x"15085776",
1866 => x"752ea338",
1867 => x"841708fc",
1868 => x"06707a31",
1869 => x"5556738f",
1870 => x"2483ca38",
1871 => x"73802584",
1872 => x"81388c17",
1873 => x"08577675",
1874 => x"2e098106",
1875 => x"df388815",
1876 => x"811b7083",
1877 => x"06555b55",
1878 => x"72c9387c",
1879 => x"83065372",
1880 => x"802efdb8",
1881 => x"38ff1df8",
1882 => x"19595d88",
1883 => x"1808782e",
1884 => x"ea38fdb5",
1885 => x"39831a53",
1886 => x"fc963983",
1887 => x"1470822c",
1888 => x"81712b80",
1889 => x"d5bc0807",
1890 => x"7080d5b8",
1891 => x"0b84050c",
1892 => x"76101010",
1893 => x"80d5b805",
1894 => x"88110859",
1895 => x"5b5e5153",
1896 => x"fee13980",
1897 => x"d4fc0817",
1898 => x"58b00876",
1899 => x"2e818d38",
1900 => x"80d5ac08",
1901 => x"ff2e83ec",
1902 => x"38737631",
1903 => x"1880d4fc",
1904 => x"0c738706",
1905 => x"70575372",
1906 => x"802e8838",
1907 => x"88733170",
1908 => x"15555676",
1909 => x"149fff06",
1910 => x"a0807131",
1911 => x"1770547f",
1912 => x"53575384",
1913 => x"e43fb008",
1914 => x"53b008ff",
1915 => x"2e81a038",
1916 => x"80d4fc08",
1917 => x"167080d4",
1918 => x"fc0c7475",
1919 => x"80d5b80b",
1920 => x"88050c74",
1921 => x"76311870",
1922 => x"81075155",
1923 => x"56587b80",
1924 => x"d5b82e83",
1925 => x"9c38798f",
1926 => x"2682cb38",
1927 => x"810b8415",
1928 => x"0c841508",
1929 => x"fc06707a",
1930 => x"317a7226",
1931 => x"8f722507",
1932 => x"52555372",
1933 => x"802efcf9",
1934 => x"3880db39",
1935 => x"b0089fff",
1936 => x"065372fe",
1937 => x"eb387780",
1938 => x"d4fc0c80",
1939 => x"d5b80b88",
1940 => x"05087b18",
1941 => x"81078412",
1942 => x"0c5580d5",
1943 => x"a8087827",
1944 => x"86387780",
1945 => x"d5a80c80",
1946 => x"d5a40878",
1947 => x"27fcac38",
1948 => x"7780d5a4",
1949 => x"0c841508",
1950 => x"fc06707a",
1951 => x"317a7226",
1952 => x"8f722507",
1953 => x"52555372",
1954 => x"802efca5",
1955 => x"38883980",
1956 => x"745456fe",
1957 => x"db397d51",
1958 => x"83ae3f80",
1959 => x"0bb00c8f",
1960 => x"3d0d0473",
1961 => x"53807424",
1962 => x"a9387282",
1963 => x"2c81712b",
1964 => x"80d5bc08",
1965 => x"077080d5",
1966 => x"b80b8405",
1967 => x"0c5d5377",
1968 => x"8c180c74",
1969 => x"88180c76",
1970 => x"88190c76",
1971 => x"8c160cf9",
1972 => x"b7398314",
1973 => x"70822c81",
1974 => x"712b80d5",
1975 => x"bc080770",
1976 => x"80d5b80b",
1977 => x"84050c5e",
1978 => x"5153d439",
1979 => x"7b7b0653",
1980 => x"72fca338",
1981 => x"841a7b10",
1982 => x"5c5af139",
1983 => x"ff1a8111",
1984 => x"515af7b9",
1985 => x"39781779",
1986 => x"81078419",
1987 => x"0c8c1808",
1988 => x"88190871",
1989 => x"8c120c88",
1990 => x"120c5970",
1991 => x"80d5cc0c",
1992 => x"7080d5c8",
1993 => x"0c80d5c0",
1994 => x"0b8c120c",
1995 => x"8c110888",
1996 => x"120c7481",
1997 => x"0784120c",
1998 => x"74117571",
1999 => x"0c5153f9",
2000 => x"bd397517",
2001 => x"84110881",
2002 => x"0784120c",
2003 => x"538c1708",
2004 => x"88180871",
2005 => x"8c120c88",
2006 => x"120c587d",
2007 => x"5181e93f",
2008 => x"881754f5",
2009 => x"cf397284",
2010 => x"150cf41a",
2011 => x"f8067084",
2012 => x"1e088106",
2013 => x"07841e0c",
2014 => x"701d545b",
2015 => x"850b8414",
2016 => x"0c850b88",
2017 => x"140c8f7b",
2018 => x"27fdcf38",
2019 => x"881c527d",
2020 => x"51ec9e3f",
2021 => x"80d5b80b",
2022 => x"88050880",
2023 => x"d4fc0859",
2024 => x"55fdb739",
2025 => x"7780d4fc",
2026 => x"0c7380d5",
2027 => x"ac0cfc91",
2028 => x"39728415",
2029 => x"0cfda339",
2030 => x"fc3d0d76",
2031 => x"7971028c",
2032 => x"059f0533",
2033 => x"57555355",
2034 => x"8372278a",
2035 => x"38748306",
2036 => x"5170802e",
2037 => x"a238ff12",
2038 => x"5271ff2e",
2039 => x"93387373",
2040 => x"70810555",
2041 => x"34ff1252",
2042 => x"71ff2e09",
2043 => x"8106ef38",
2044 => x"74b00c86",
2045 => x"3d0d0474",
2046 => x"74882b75",
2047 => x"07707190",
2048 => x"2b075154",
2049 => x"518f7227",
2050 => x"a5387271",
2051 => x"70840553",
2052 => x"0c727170",
2053 => x"8405530c",
2054 => x"72717084",
2055 => x"05530c72",
2056 => x"71708405",
2057 => x"530cf012",
2058 => x"52718f26",
2059 => x"dd388372",
2060 => x"27903872",
2061 => x"71708405",
2062 => x"530cfc12",
2063 => x"52718326",
2064 => x"f2387053",
2065 => x"ff903904",
2066 => x"04fd3d0d",
2067 => x"800b80dd",
2068 => x"f40c7651",
2069 => x"84ee3fb0",
2070 => x"0853b008",
2071 => x"ff2e8838",
2072 => x"72b00c85",
2073 => x"3d0d0480",
2074 => x"ddf40854",
2075 => x"73802ef0",
2076 => x"38757471",
2077 => x"0c5272b0",
2078 => x"0c853d0d",
2079 => x"04f93d0d",
2080 => x"797c557b",
2081 => x"548e1122",
2082 => x"70902b70",
2083 => x"902c5557",
2084 => x"80cdfc08",
2085 => x"53585683",
2086 => x"f33fb008",
2087 => x"57800bb0",
2088 => x"08249338",
2089 => x"80d01608",
2090 => x"b0080580",
2091 => x"d0170c76",
2092 => x"b00c893d",
2093 => x"0d048c16",
2094 => x"2283dfff",
2095 => x"0655748c",
2096 => x"172376b0",
2097 => x"0c893d0d",
2098 => x"04fa3d0d",
2099 => x"788c1122",
2100 => x"70882a70",
2101 => x"81065157",
2102 => x"585674a9",
2103 => x"388c1622",
2104 => x"83dfff06",
2105 => x"55748c17",
2106 => x"237a5479",
2107 => x"538e1622",
2108 => x"70902b70",
2109 => x"902c5456",
2110 => x"80cdfc08",
2111 => x"525681b2",
2112 => x"3f883d0d",
2113 => x"04825480",
2114 => x"538e1622",
2115 => x"70902b70",
2116 => x"902c5456",
2117 => x"80cdfc08",
2118 => x"525782b8",
2119 => x"3f8c1622",
2120 => x"83dfff06",
2121 => x"55748c17",
2122 => x"237a5479",
2123 => x"538e1622",
2124 => x"70902b70",
2125 => x"902c5456",
2126 => x"80cdfc08",
2127 => x"525680f2",
2128 => x"3f883d0d",
2129 => x"04f93d0d",
2130 => x"797c557b",
2131 => x"548e1122",
2132 => x"70902b70",
2133 => x"902c5557",
2134 => x"80cdfc08",
2135 => x"53585681",
2136 => x"f33fb008",
2137 => x"57b008ff",
2138 => x"2e99388c",
2139 => x"1622a080",
2140 => x"0755748c",
2141 => x"1723b008",
2142 => x"80d0170c",
2143 => x"76b00c89",
2144 => x"3d0d048c",
2145 => x"162283df",
2146 => x"ff065574",
2147 => x"8c172376",
2148 => x"b00c893d",
2149 => x"0d04fe3d",
2150 => x"0d748e11",
2151 => x"2270902b",
2152 => x"70902c55",
2153 => x"51515380",
2154 => x"cdfc0851",
2155 => x"bd3f843d",
2156 => x"0d04fb3d",
2157 => x"0d800b80",
2158 => x"ddf40c7a",
2159 => x"53795278",
2160 => x"5182f93f",
2161 => x"b00855b0",
2162 => x"08ff2e88",
2163 => x"3874b00c",
2164 => x"873d0d04",
2165 => x"80ddf408",
2166 => x"5675802e",
2167 => x"f0387776",
2168 => x"710c5474",
2169 => x"b00c873d",
2170 => x"0d04fd3d",
2171 => x"0d800b80",
2172 => x"ddf40c76",
2173 => x"5184c33f",
2174 => x"b00853b0",
2175 => x"08ff2e88",
2176 => x"3872b00c",
2177 => x"853d0d04",
2178 => x"80ddf408",
2179 => x"5473802e",
2180 => x"f0387574",
2181 => x"710c5272",
2182 => x"b00c853d",
2183 => x"0d04fc3d",
2184 => x"0d800b80",
2185 => x"ddf40c78",
2186 => x"52775186",
2187 => x"ab3fb008",
2188 => x"54b008ff",
2189 => x"2e883873",
2190 => x"b00c863d",
2191 => x"0d0480dd",
2192 => x"f4085574",
2193 => x"802ef038",
2194 => x"7675710c",
2195 => x"5373b00c",
2196 => x"863d0d04",
2197 => x"fb3d0d80",
2198 => x"0b80ddf4",
2199 => x"0c7a5379",
2200 => x"52785184",
2201 => x"873fb008",
2202 => x"55b008ff",
2203 => x"2e883874",
2204 => x"b00c873d",
2205 => x"0d0480dd",
2206 => x"f4085675",
2207 => x"802ef038",
2208 => x"7776710c",
2209 => x"5474b00c",
2210 => x"873d0d04",
2211 => x"fb3d0d80",
2212 => x"0b80ddf4",
2213 => x"0c7a5379",
2214 => x"52785182",
2215 => x"933fb008",
2216 => x"55b008ff",
2217 => x"2e883874",
2218 => x"b00c873d",
2219 => x"0d0480dd",
2220 => x"f4085675",
2221 => x"802ef038",
2222 => x"7776710c",
2223 => x"5474b00c",
2224 => x"873d0d04",
2225 => x"fe3d0d80",
2226 => x"dde80851",
2227 => x"708a3880",
2228 => x"ddf87080",
2229 => x"dde80c51",
2230 => x"70751252",
2231 => x"52ff5370",
2232 => x"87fb8080",
2233 => x"26883870",
2234 => x"80dde80c",
2235 => x"715372b0",
2236 => x"0c843d0d",
2237 => x"04fd3d0d",
2238 => x"800b80cd",
2239 => x"f0085454",
2240 => x"72812e9b",
2241 => x"387380dd",
2242 => x"ec0cc3da",
2243 => x"3fc1f13f",
2244 => x"80ddc052",
2245 => x"8151c5b0",
2246 => x"3fb00851",
2247 => x"85ba3f72",
2248 => x"80ddec0c",
2249 => x"c3c03fc1",
2250 => x"d73f80dd",
2251 => x"c0528151",
2252 => x"c5963fb0",
2253 => x"085185a0",
2254 => x"3f00ff39",
2255 => x"f53d0d7e",
2256 => x"6080ddec",
2257 => x"08705b58",
2258 => x"5b5b7580",
2259 => x"c238777a",
2260 => x"25a13877",
2261 => x"1b703370",
2262 => x"81ff0658",
2263 => x"5859758a",
2264 => x"2e983876",
2265 => x"81ff0651",
2266 => x"c2db3f81",
2267 => x"18587978",
2268 => x"24e13879",
2269 => x"b00c8d3d",
2270 => x"0d048d51",
2271 => x"c2c73f78",
2272 => x"337081ff",
2273 => x"065257c2",
2274 => x"bc3f8118",
2275 => x"58e03979",
2276 => x"557a547d",
2277 => x"5385528d",
2278 => x"3dfc0551",
2279 => x"c1a43fb0",
2280 => x"085684ad",
2281 => x"3f7bb008",
2282 => x"0c75b00c",
2283 => x"8d3d0d04",
2284 => x"f63d0d7d",
2285 => x"7f80ddec",
2286 => x"08705b58",
2287 => x"5a5a7580",
2288 => x"c1387779",
2289 => x"25b338c1",
2290 => x"d73fb008",
2291 => x"81ff0670",
2292 => x"8d327030",
2293 => x"709f2a51",
2294 => x"51575776",
2295 => x"8a2e80c3",
2296 => x"3875802e",
2297 => x"be38771a",
2298 => x"56767634",
2299 => x"7651c1d5",
2300 => x"3f811858",
2301 => x"787824cf",
2302 => x"38775675",
2303 => x"b00c8c3d",
2304 => x"0d047855",
2305 => x"79547c53",
2306 => x"84528c3d",
2307 => x"fc0551c0",
2308 => x"b13fb008",
2309 => x"5683ba3f",
2310 => x"7ab0080c",
2311 => x"75b00c8c",
2312 => x"3d0d0477",
2313 => x"1a568a76",
2314 => x"34811858",
2315 => x"8d51c195",
2316 => x"3f8a51c1",
2317 => x"903f7756",
2318 => x"c239fb3d",
2319 => x"0d80ddec",
2320 => x"08705654",
2321 => x"73883874",
2322 => x"b00c873d",
2323 => x"0d047753",
2324 => x"8352873d",
2325 => x"fc0551ff",
2326 => x"bfe83fb0",
2327 => x"085482f1",
2328 => x"3f75b008",
2329 => x"0c73b00c",
2330 => x"873d0d04",
2331 => x"fa3d0d80",
2332 => x"ddec0880",
2333 => x"2ea3387a",
2334 => x"55795478",
2335 => x"53865288",
2336 => x"3dfc0551",
2337 => x"ffbfbb3f",
2338 => x"b0085682",
2339 => x"c43f76b0",
2340 => x"080c75b0",
2341 => x"0c883d0d",
2342 => x"0482b63f",
2343 => x"9d0bb008",
2344 => x"0cff0bb0",
2345 => x"0c883d0d",
2346 => x"04fb3d0d",
2347 => x"77795656",
2348 => x"80705454",
2349 => x"7375259f",
2350 => x"38741010",
2351 => x"10f80552",
2352 => x"72167033",
2353 => x"70742b76",
2354 => x"078116f8",
2355 => x"16565656",
2356 => x"51517473",
2357 => x"24ea3873",
2358 => x"b00c873d",
2359 => x"0d04fc3d",
2360 => x"0d767855",
2361 => x"55bc5380",
2362 => x"527351f5",
2363 => x"cb3f8452",
2364 => x"7451ffb5",
2365 => x"3fb00874",
2366 => x"23845284",
2367 => x"1551ffa9",
2368 => x"3fb00882",
2369 => x"15238452",
2370 => x"881551ff",
2371 => x"9c3fb008",
2372 => x"84150c84",
2373 => x"528c1551",
2374 => x"ff8f3fb0",
2375 => x"08881523",
2376 => x"84529015",
2377 => x"51ff823f",
2378 => x"b0088a15",
2379 => x"23845294",
2380 => x"1551fef5",
2381 => x"3fb0088c",
2382 => x"15238452",
2383 => x"981551fe",
2384 => x"e83fb008",
2385 => x"8e152388",
2386 => x"529c1551",
2387 => x"fedb3fb0",
2388 => x"0890150c",
2389 => x"863d0d04",
2390 => x"e93d0d6a",
2391 => x"80ddec08",
2392 => x"57577593",
2393 => x"3880c080",
2394 => x"0b84180c",
2395 => x"75ac180c",
2396 => x"75b00c99",
2397 => x"3d0d0489",
2398 => x"3d70556a",
2399 => x"54558a52",
2400 => x"993dffbc",
2401 => x"0551ffbd",
2402 => x"b93fb008",
2403 => x"77537552",
2404 => x"56fecb3f",
2405 => x"bc3f77b0",
2406 => x"080c75b0",
2407 => x"0c993d0d",
2408 => x"04fc3d0d",
2409 => x"815480dd",
2410 => x"ec088838",
2411 => x"73b00c86",
2412 => x"3d0d0476",
2413 => x"5397b952",
2414 => x"863dfc05",
2415 => x"51ffbd82",
2416 => x"3fb00854",
2417 => x"8c3f74b0",
2418 => x"080c73b0",
2419 => x"0c863d0d",
2420 => x"0480cdfc",
2421 => x"08b00c04",
2422 => x"f73d0d7b",
2423 => x"80cdfc08",
2424 => x"82c81108",
2425 => x"5a545a77",
2426 => x"802e80da",
2427 => x"38818818",
2428 => x"841908ff",
2429 => x"0581712b",
2430 => x"59555980",
2431 => x"742480ea",
2432 => x"38807424",
2433 => x"b5387382",
2434 => x"2b781188",
2435 => x"05565681",
2436 => x"80190877",
2437 => x"06537280",
2438 => x"2eb63878",
2439 => x"16700853",
2440 => x"53795174",
2441 => x"0853722d",
2442 => x"ff14fc17",
2443 => x"fc177981",
2444 => x"2c5a5757",
2445 => x"54738025",
2446 => x"d6387708",
2447 => x"5877ffad",
2448 => x"3880cdfc",
2449 => x"0853bc13",
2450 => x"08a53879",
2451 => x"51f9ea3f",
2452 => x"74085372",
2453 => x"2dff14fc",
2454 => x"17fc1779",
2455 => x"812c5a57",
2456 => x"57547380",
2457 => x"25ffa838",
2458 => x"d1398057",
2459 => x"ff933972",
2460 => x"51bc1308",
2461 => x"53722d79",
2462 => x"51f9be3f",
2463 => x"ff3d0d80",
2464 => x"ddc80bfc",
2465 => x"05700852",
2466 => x"5270ff2e",
2467 => x"9138702d",
2468 => x"fc127008",
2469 => x"525270ff",
2470 => x"2e098106",
2471 => x"f138833d",
2472 => x"0d0404ff",
2473 => x"bdab3f04",
2474 => x"00ffffff",
2475 => x"ff00ffff",
2476 => x"ffff00ff",
2477 => x"ffffff00",
2478 => x"00000040",
2479 => x"476f7420",
2480 => x"696e7465",
2481 => x"72727570",
2482 => x"740a0000",
2483 => x"4e6f2069",
2484 => x"6e746572",
2485 => x"72757074",
2486 => x"0a000000",
2487 => x"43000000",
2488 => x"64756d6d",
2489 => x"792e6578",
2490 => x"65000000",
2491 => x"00000000",
2492 => x"00000000",
2493 => x"00000000",
2494 => x"00002ed0",
2495 => x"00002700",
2496 => x"00000000",
2497 => x"00002968",
2498 => x"000029c4",
2499 => x"00002a20",
2500 => x"00000000",
2501 => x"00000000",
2502 => x"00000000",
2503 => x"00000000",
2504 => x"00000000",
2505 => x"00000000",
2506 => x"00000000",
2507 => x"00000000",
2508 => x"00000000",
2509 => x"000026dc",
2510 => x"00000000",
2511 => x"00000000",
2512 => x"00000000",
2513 => x"00000000",
2514 => x"00000000",
2515 => x"00000000",
2516 => x"00000000",
2517 => x"00000000",
2518 => x"00000000",
2519 => x"00000000",
2520 => x"00000000",
2521 => x"00000000",
2522 => x"00000000",
2523 => x"00000000",
2524 => x"00000000",
2525 => x"00000000",
2526 => x"00000000",
2527 => x"00000000",
2528 => x"00000000",
2529 => x"00000000",
2530 => x"00000000",
2531 => x"00000000",
2532 => x"00000000",
2533 => x"00000000",
2534 => x"00000000",
2535 => x"00000000",
2536 => x"00000000",
2537 => x"00000000",
2538 => x"00000001",
2539 => x"330eabcd",
2540 => x"1234e66d",
2541 => x"deec0005",
2542 => x"000b0000",
2543 => x"00000000",
2544 => x"00000000",
2545 => x"00000000",
2546 => x"00000000",
2547 => x"00000000",
2548 => x"00000000",
2549 => x"00000000",
2550 => x"00000000",
2551 => x"00000000",
2552 => x"00000000",
2553 => x"00000000",
2554 => x"00000000",
2555 => x"00000000",
2556 => x"00000000",
2557 => x"00000000",
2558 => x"00000000",
2559 => x"00000000",
2560 => x"00000000",
2561 => x"00000000",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"00000000",
2568 => x"00000000",
2569 => x"00000000",
2570 => x"00000000",
2571 => x"00000000",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000000",
2586 => x"00000000",
2587 => x"00000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000000",
2597 => x"00000000",
2598 => x"00000000",
2599 => x"00000000",
2600 => x"00000000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"ffffffff",
2732 => x"00000000",
2733 => x"00020000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00002ab8",
2737 => x"00002ab8",
2738 => x"00002ac0",
2739 => x"00002ac0",
2740 => x"00002ac8",
2741 => x"00002ac8",
2742 => x"00002ad0",
2743 => x"00002ad0",
2744 => x"00002ad8",
2745 => x"00002ad8",
2746 => x"00002ae0",
2747 => x"00002ae0",
2748 => x"00002ae8",
2749 => x"00002ae8",
2750 => x"00002af0",
2751 => x"00002af0",
2752 => x"00002af8",
2753 => x"00002af8",
2754 => x"00002b00",
2755 => x"00002b00",
2756 => x"00002b08",
2757 => x"00002b08",
2758 => x"00002b10",
2759 => x"00002b10",
2760 => x"00002b18",
2761 => x"00002b18",
2762 => x"00002b20",
2763 => x"00002b20",
2764 => x"00002b28",
2765 => x"00002b28",
2766 => x"00002b30",
2767 => x"00002b30",
2768 => x"00002b38",
2769 => x"00002b38",
2770 => x"00002b40",
2771 => x"00002b40",
2772 => x"00002b48",
2773 => x"00002b48",
2774 => x"00002b50",
2775 => x"00002b50",
2776 => x"00002b58",
2777 => x"00002b58",
2778 => x"00002b60",
2779 => x"00002b60",
2780 => x"00002b68",
2781 => x"00002b68",
2782 => x"00002b70",
2783 => x"00002b70",
2784 => x"00002b78",
2785 => x"00002b78",
2786 => x"00002b80",
2787 => x"00002b80",
2788 => x"00002b88",
2789 => x"00002b88",
2790 => x"00002b90",
2791 => x"00002b90",
2792 => x"00002b98",
2793 => x"00002b98",
2794 => x"00002ba0",
2795 => x"00002ba0",
2796 => x"00002ba8",
2797 => x"00002ba8",
2798 => x"00002bb0",
2799 => x"00002bb0",
2800 => x"00002bb8",
2801 => x"00002bb8",
2802 => x"00002bc0",
2803 => x"00002bc0",
2804 => x"00002bc8",
2805 => x"00002bc8",
2806 => x"00002bd0",
2807 => x"00002bd0",
2808 => x"00002bd8",
2809 => x"00002bd8",
2810 => x"00002be0",
2811 => x"00002be0",
2812 => x"00002be8",
2813 => x"00002be8",
2814 => x"00002bf0",
2815 => x"00002bf0",
2816 => x"00002bf8",
2817 => x"00002bf8",
2818 => x"00002c00",
2819 => x"00002c00",
2820 => x"00002c08",
2821 => x"00002c08",
2822 => x"00002c10",
2823 => x"00002c10",
2824 => x"00002c18",
2825 => x"00002c18",
2826 => x"00002c20",
2827 => x"00002c20",
2828 => x"00002c28",
2829 => x"00002c28",
2830 => x"00002c30",
2831 => x"00002c30",
2832 => x"00002c38",
2833 => x"00002c38",
2834 => x"00002c40",
2835 => x"00002c40",
2836 => x"00002c48",
2837 => x"00002c48",
2838 => x"00002c50",
2839 => x"00002c50",
2840 => x"00002c58",
2841 => x"00002c58",
2842 => x"00002c60",
2843 => x"00002c60",
2844 => x"00002c68",
2845 => x"00002c68",
2846 => x"00002c70",
2847 => x"00002c70",
2848 => x"00002c78",
2849 => x"00002c78",
2850 => x"00002c80",
2851 => x"00002c80",
2852 => x"00002c88",
2853 => x"00002c88",
2854 => x"00002c90",
2855 => x"00002c90",
2856 => x"00002c98",
2857 => x"00002c98",
2858 => x"00002ca0",
2859 => x"00002ca0",
2860 => x"00002ca8",
2861 => x"00002ca8",
2862 => x"00002cb0",
2863 => x"00002cb0",
2864 => x"00002cb8",
2865 => x"00002cb8",
2866 => x"00002cc0",
2867 => x"00002cc0",
2868 => x"00002cc8",
2869 => x"00002cc8",
2870 => x"00002cd0",
2871 => x"00002cd0",
2872 => x"00002cd8",
2873 => x"00002cd8",
2874 => x"00002ce0",
2875 => x"00002ce0",
2876 => x"00002ce8",
2877 => x"00002ce8",
2878 => x"00002cf0",
2879 => x"00002cf0",
2880 => x"00002cf8",
2881 => x"00002cf8",
2882 => x"00002d00",
2883 => x"00002d00",
2884 => x"00002d08",
2885 => x"00002d08",
2886 => x"00002d10",
2887 => x"00002d10",
2888 => x"00002d18",
2889 => x"00002d18",
2890 => x"00002d20",
2891 => x"00002d20",
2892 => x"00002d28",
2893 => x"00002d28",
2894 => x"00002d30",
2895 => x"00002d30",
2896 => x"00002d38",
2897 => x"00002d38",
2898 => x"00002d40",
2899 => x"00002d40",
2900 => x"00002d48",
2901 => x"00002d48",
2902 => x"00002d50",
2903 => x"00002d50",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"000026e0",
2993 => x"ffffffff",
2994 => x"00000000",
2995 => x"ffffffff",
2996 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

