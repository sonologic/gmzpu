------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80d0f40c",
3 => x"3a0b0b80",
4 => x"c8d00400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d0",
162 => x"90738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d0f00c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c7de3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8ffe2d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8ecc2d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80e0e0",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80e0",
307 => x"e0085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480d0",
314 => x"f008802e",
315 => x"a43880d0",
316 => x"f408822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80e0e00c",
320 => x"82a0800b",
321 => x"80e0e40c",
322 => x"8290800b",
323 => x"80e0e80c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80e0e0",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"e0e40cf8",
330 => x"80808480",
331 => x"0b80e0e8",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80e0",
335 => x"e00c80c0",
336 => x"a880940b",
337 => x"80e0e40c",
338 => x"80d0a00b",
339 => x"80e0e80c",
340 => x"04ff3d0d",
341 => x"80e0ec33",
342 => x"5170a738",
343 => x"80d0fc08",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"d0fc0c70",
348 => x"2d80d0fc",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80e0",
352 => x"ec34833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80e0dc08",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"e0dc510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404803d",
366 => x"0d80e0f8",
367 => x"08811180",
368 => x"e0f80c51",
369 => x"823d0d04",
370 => x"f73d0d7b",
371 => x"54870b89",
372 => x"3d80d180",
373 => x"08585855",
374 => x"7417748f",
375 => x"06175353",
376 => x"71337334",
377 => x"73842aff",
378 => x"16565474",
379 => x"8025e938",
380 => x"800b8b3d",
381 => x"34765188",
382 => x"aa3f8b3d",
383 => x"0d04e93d",
384 => x"0d80e0f8",
385 => x"08973d95",
386 => x"3d933d91",
387 => x"3d80e0f8",
388 => x"08575c5c",
389 => x"5c5c5c7b",
390 => x"722e828b",
391 => x"3880d0b8",
392 => x"5188803f",
393 => x"80e0f808",
394 => x"8c808008",
395 => x"8c808408",
396 => x"80d0c854",
397 => x"59545c87",
398 => x"ea3f7254",
399 => x"870b80d1",
400 => x"80085755",
401 => x"741b748f",
402 => x"06175353",
403 => x"71337334",
404 => x"73842aff",
405 => x"16565474",
406 => x"8025e938",
407 => x"800b993d",
408 => x"347a5187",
409 => x"be3f80d0",
410 => x"cc5187b7",
411 => x"3f765487",
412 => x"0b80d180",
413 => x"08575574",
414 => x"1a748f06",
415 => x"17545772",
416 => x"33773473",
417 => x"842aff16",
418 => x"56547480",
419 => x"25e93880",
420 => x"0b963d34",
421 => x"7951878b",
422 => x"3f800b8c",
423 => x"80800c81",
424 => x"91d1acf8",
425 => x"0b8c8084",
426 => x"0c8c8080",
427 => x"088c8084",
428 => x"0880d0c8",
429 => x"53585586",
430 => x"ea3f7454",
431 => x"870b80d1",
432 => x"80085755",
433 => x"7419748f",
434 => x"06175353",
435 => x"71337334",
436 => x"73842aff",
437 => x"16565474",
438 => x"8025e938",
439 => x"800b933d",
440 => x"34785186",
441 => x"be3f80d0",
442 => x"cc5186b7",
443 => x"3f765487",
444 => x"0b80d180",
445 => x"08575574",
446 => x"18748f06",
447 => x"17545772",
448 => x"33773473",
449 => x"842aff16",
450 => x"56547480",
451 => x"25e93880",
452 => x"0b903d34",
453 => x"7751868b",
454 => x"3f80e0f8",
455 => x"08527b72",
456 => x"2e098106",
457 => x"fdf73880",
458 => x"d0d05185",
459 => x"f63f8c80",
460 => x"80088c80",
461 => x"840880d0",
462 => x"c8535853",
463 => x"85e53f72",
464 => x"54870b80",
465 => x"d1800857",
466 => x"55fdf939",
467 => x"bc0802bc",
468 => x"0cf93d0d",
469 => x"800bbc08",
470 => x"fc050cbc",
471 => x"08880508",
472 => x"8025ab38",
473 => x"bc088805",
474 => x"0830bc08",
475 => x"88050c80",
476 => x"0bbc08f4",
477 => x"050cbc08",
478 => x"fc050888",
479 => x"38810bbc",
480 => x"08f4050c",
481 => x"bc08f405",
482 => x"08bc08fc",
483 => x"050cbc08",
484 => x"8c050880",
485 => x"25ab38bc",
486 => x"088c0508",
487 => x"30bc088c",
488 => x"050c800b",
489 => x"bc08f005",
490 => x"0cbc08fc",
491 => x"05088838",
492 => x"810bbc08",
493 => x"f0050cbc",
494 => x"08f00508",
495 => x"bc08fc05",
496 => x"0c8053bc",
497 => x"088c0508",
498 => x"52bc0888",
499 => x"05085181",
500 => x"a73fb008",
501 => x"70bc08f8",
502 => x"050c54bc",
503 => x"08fc0508",
504 => x"802e8c38",
505 => x"bc08f805",
506 => x"0830bc08",
507 => x"f8050cbc",
508 => x"08f80508",
509 => x"70b00c54",
510 => x"893d0dbc",
511 => x"0c04bc08",
512 => x"02bc0cfb",
513 => x"3d0d800b",
514 => x"bc08fc05",
515 => x"0cbc0888",
516 => x"05088025",
517 => x"9338bc08",
518 => x"88050830",
519 => x"bc088805",
520 => x"0c810bbc",
521 => x"08fc050c",
522 => x"bc088c05",
523 => x"0880258c",
524 => x"38bc088c",
525 => x"050830bc",
526 => x"088c050c",
527 => x"8153bc08",
528 => x"8c050852",
529 => x"bc088805",
530 => x"0851ad3f",
531 => x"b00870bc",
532 => x"08f8050c",
533 => x"54bc08fc",
534 => x"0508802e",
535 => x"8c38bc08",
536 => x"f8050830",
537 => x"bc08f805",
538 => x"0cbc08f8",
539 => x"050870b0",
540 => x"0c54873d",
541 => x"0dbc0c04",
542 => x"bc0802bc",
543 => x"0cfd3d0d",
544 => x"810bbc08",
545 => x"fc050c80",
546 => x"0bbc08f8",
547 => x"050cbc08",
548 => x"8c0508bc",
549 => x"08880508",
550 => x"27ac38bc",
551 => x"08fc0508",
552 => x"802ea338",
553 => x"800bbc08",
554 => x"8c050824",
555 => x"9938bc08",
556 => x"8c050810",
557 => x"bc088c05",
558 => x"0cbc08fc",
559 => x"050810bc",
560 => x"08fc050c",
561 => x"c939bc08",
562 => x"fc050880",
563 => x"2e80c938",
564 => x"bc088c05",
565 => x"08bc0888",
566 => x"050826a1",
567 => x"38bc0888",
568 => x"0508bc08",
569 => x"8c050831",
570 => x"bc088805",
571 => x"0cbc08f8",
572 => x"0508bc08",
573 => x"fc050807",
574 => x"bc08f805",
575 => x"0cbc08fc",
576 => x"0508812a",
577 => x"bc08fc05",
578 => x"0cbc088c",
579 => x"0508812a",
580 => x"bc088c05",
581 => x"0cffaf39",
582 => x"bc089005",
583 => x"08802e8f",
584 => x"38bc0888",
585 => x"050870bc",
586 => x"08f4050c",
587 => x"518d39bc",
588 => x"08f80508",
589 => x"70bc08f4",
590 => x"050c51bc",
591 => x"08f40508",
592 => x"b00c853d",
593 => x"0dbc0c04",
594 => x"fc3d0d76",
595 => x"70797b55",
596 => x"5555558f",
597 => x"72278c38",
598 => x"72750783",
599 => x"06517080",
600 => x"2ea738ff",
601 => x"125271ff",
602 => x"2e983872",
603 => x"70810554",
604 => x"33747081",
605 => x"055634ff",
606 => x"125271ff",
607 => x"2e098106",
608 => x"ea3874b0",
609 => x"0c863d0d",
610 => x"04745172",
611 => x"70840554",
612 => x"08717084",
613 => x"05530c72",
614 => x"70840554",
615 => x"08717084",
616 => x"05530c72",
617 => x"70840554",
618 => x"08717084",
619 => x"05530c72",
620 => x"70840554",
621 => x"08717084",
622 => x"05530cf0",
623 => x"1252718f",
624 => x"26c93883",
625 => x"72279538",
626 => x"72708405",
627 => x"54087170",
628 => x"8405530c",
629 => x"fc125271",
630 => x"8326ed38",
631 => x"7054ff83",
632 => x"39f73d0d",
633 => x"7c705253",
634 => x"80ca3f72",
635 => x"54b00855",
636 => x"0b0b80d0",
637 => x"dc568157",
638 => x"b0088105",
639 => x"5a8b3de4",
640 => x"11595382",
641 => x"59f41352",
642 => x"7b881108",
643 => x"52538183",
644 => x"3fb00830",
645 => x"70b00807",
646 => x"9f2c8a07",
647 => x"b00c538b",
648 => x"3d0d04ff",
649 => x"3d0d7352",
650 => x"80d18408",
651 => x"51ffb23f",
652 => x"833d0d04",
653 => x"fd3d0d75",
654 => x"70718306",
655 => x"53555270",
656 => x"b8387170",
657 => x"087009f7",
658 => x"fbfdff12",
659 => x"0670f884",
660 => x"82818006",
661 => x"51515253",
662 => x"709d3884",
663 => x"13700870",
664 => x"09f7fbfd",
665 => x"ff120670",
666 => x"f8848281",
667 => x"80065151",
668 => x"52537080",
669 => x"2ee53872",
670 => x"52713351",
671 => x"70802e8a",
672 => x"38811270",
673 => x"33525270",
674 => x"f8387174",
675 => x"31b00c85",
676 => x"3d0d04f2",
677 => x"3d0d6062",
678 => x"88110870",
679 => x"57575f5a",
680 => x"74802e81",
681 => x"8f388c1a",
682 => x"2270832a",
683 => x"81327081",
684 => x"06515558",
685 => x"73863890",
686 => x"1a089138",
687 => x"795190a1",
688 => x"3fff54b0",
689 => x"0880ed38",
690 => x"8c1a2258",
691 => x"7d085780",
692 => x"7883ffff",
693 => x"0670812a",
694 => x"70810651",
695 => x"56575573",
696 => x"752e80d7",
697 => x"38749038",
698 => x"76088418",
699 => x"08881959",
700 => x"56597480",
701 => x"2ef23874",
702 => x"54888075",
703 => x"27843888",
704 => x"80547353",
705 => x"78529c1a",
706 => x"0851a41a",
707 => x"0854732d",
708 => x"800bb008",
709 => x"2582e638",
710 => x"b0081975",
711 => x"b008317f",
712 => x"880508b0",
713 => x"08317061",
714 => x"88050c56",
715 => x"565973ff",
716 => x"b4388054",
717 => x"73b00c90",
718 => x"3d0d0475",
719 => x"81327081",
720 => x"06764151",
721 => x"5473802e",
722 => x"81c13874",
723 => x"90387608",
724 => x"84180888",
725 => x"19595659",
726 => x"74802ef2",
727 => x"38881a08",
728 => x"7883ffff",
729 => x"0670892a",
730 => x"70810651",
731 => x"56595673",
732 => x"802e82fa",
733 => x"38757527",
734 => x"8d387787",
735 => x"2a708106",
736 => x"51547382",
737 => x"b5387476",
738 => x"27833874",
739 => x"56755378",
740 => x"52790851",
741 => x"85823f88",
742 => x"1a087631",
743 => x"881b0c79",
744 => x"08167a0c",
745 => x"74567519",
746 => x"7577317f",
747 => x"88050878",
748 => x"31706188",
749 => x"050c5656",
750 => x"5973802e",
751 => x"fef4388c",
752 => x"1a2258ff",
753 => x"86397778",
754 => x"5479537b",
755 => x"525684c8",
756 => x"3f881a08",
757 => x"7831881b",
758 => x"0c790818",
759 => x"7a0c7c76",
760 => x"315d7c8e",
761 => x"3879518f",
762 => x"db3fb008",
763 => x"818f38b0",
764 => x"085f7519",
765 => x"7577317f",
766 => x"88050878",
767 => x"31706188",
768 => x"050c5656",
769 => x"5973802e",
770 => x"fea83874",
771 => x"81833876",
772 => x"08841808",
773 => x"88195956",
774 => x"5974802e",
775 => x"f2387453",
776 => x"8a527851",
777 => x"82d33fb0",
778 => x"08793181",
779 => x"055db008",
780 => x"84388115",
781 => x"5d815f7c",
782 => x"58747d27",
783 => x"83387458",
784 => x"941a0888",
785 => x"1b081157",
786 => x"5c807a08",
787 => x"5c54901a",
788 => x"087b2783",
789 => x"38815475",
790 => x"78258438",
791 => x"73ba387b",
792 => x"7824fee2",
793 => x"387b5378",
794 => x"529c1a08",
795 => x"51a41a08",
796 => x"54732db0",
797 => x"0856b008",
798 => x"8024fee2",
799 => x"388c1a22",
800 => x"80c00754",
801 => x"738c1b23",
802 => x"ff5473b0",
803 => x"0c903d0d",
804 => x"047effa3",
805 => x"38ff8739",
806 => x"75537852",
807 => x"7a5182f8",
808 => x"3f790816",
809 => x"7a0c7951",
810 => x"8e9a3fb0",
811 => x"08cf387c",
812 => x"76315d7c",
813 => x"febc38fe",
814 => x"ac39901a",
815 => x"087a0871",
816 => x"31761170",
817 => x"565a5752",
818 => x"80d18408",
819 => x"51848c3f",
820 => x"b008802e",
821 => x"ffa738b0",
822 => x"08901b0c",
823 => x"b008167a",
824 => x"0c77941b",
825 => x"0c74881b",
826 => x"0c7456fd",
827 => x"99397908",
828 => x"58901a08",
829 => x"78278338",
830 => x"81547575",
831 => x"27843873",
832 => x"b338941a",
833 => x"08567575",
834 => x"2680d338",
835 => x"75537852",
836 => x"9c1a0851",
837 => x"a41a0854",
838 => x"732db008",
839 => x"56b00880",
840 => x"24fd8338",
841 => x"8c1a2280",
842 => x"c0075473",
843 => x"8c1b23ff",
844 => x"54fed739",
845 => x"75537852",
846 => x"775181dc",
847 => x"3f790816",
848 => x"7a0c7951",
849 => x"8cfe3fb0",
850 => x"08802efc",
851 => x"d9388c1a",
852 => x"2280c007",
853 => x"54738c1b",
854 => x"23ff54fe",
855 => x"ad397475",
856 => x"54795378",
857 => x"525681b0",
858 => x"3f881a08",
859 => x"7531881b",
860 => x"0c790815",
861 => x"7a0cfcae",
862 => x"39fa3d0d",
863 => x"7a790288",
864 => x"05a70533",
865 => x"56525383",
866 => x"73278a38",
867 => x"70830652",
868 => x"71802ea8",
869 => x"38ff1353",
870 => x"72ff2e97",
871 => x"38703352",
872 => x"73722e91",
873 => x"388111ff",
874 => x"14545172",
875 => x"ff2e0981",
876 => x"06eb3880",
877 => x"5170b00c",
878 => x"883d0d04",
879 => x"70725755",
880 => x"83517582",
881 => x"802914ff",
882 => x"12525670",
883 => x"8025f338",
884 => x"837327bf",
885 => x"38740876",
886 => x"327009f7",
887 => x"fbfdff12",
888 => x"0670f884",
889 => x"82818006",
890 => x"51515170",
891 => x"802e9938",
892 => x"74518052",
893 => x"70335773",
894 => x"772effb9",
895 => x"38811181",
896 => x"13535183",
897 => x"7227ed38",
898 => x"fc138416",
899 => x"56537283",
900 => x"26c33874",
901 => x"51fefe39",
902 => x"fa3d0d78",
903 => x"7a7c7272",
904 => x"72575757",
905 => x"59565674",
906 => x"7627b238",
907 => x"76155175",
908 => x"7127aa38",
909 => x"707717ff",
910 => x"14545553",
911 => x"71ff2e96",
912 => x"38ff14ff",
913 => x"14545472",
914 => x"337434ff",
915 => x"125271ff",
916 => x"2e098106",
917 => x"ec3875b0",
918 => x"0c883d0d",
919 => x"04768f26",
920 => x"9738ff12",
921 => x"5271ff2e",
922 => x"ed387270",
923 => x"81055433",
924 => x"74708105",
925 => x"5634eb39",
926 => x"74760783",
927 => x"065170e2",
928 => x"38757554",
929 => x"51727084",
930 => x"05540871",
931 => x"70840553",
932 => x"0c727084",
933 => x"05540871",
934 => x"70840553",
935 => x"0c727084",
936 => x"05540871",
937 => x"70840553",
938 => x"0c727084",
939 => x"05540871",
940 => x"70840553",
941 => x"0cf01252",
942 => x"718f26c9",
943 => x"38837227",
944 => x"95387270",
945 => x"84055408",
946 => x"71708405",
947 => x"530cfc12",
948 => x"52718326",
949 => x"ed387054",
950 => x"ff8839ef",
951 => x"3d0d6365",
952 => x"67405d42",
953 => x"7b802e84",
954 => x"fa386151",
955 => x"a5b43ff8",
956 => x"1c708412",
957 => x"0870fc06",
958 => x"70628b05",
959 => x"70f80641",
960 => x"59455b5c",
961 => x"41579674",
962 => x"2782c338",
963 => x"807b247e",
964 => x"7c260759",
965 => x"80547874",
966 => x"2e098106",
967 => x"82a93877",
968 => x"7b2581fc",
969 => x"38771780",
970 => x"d8c00b88",
971 => x"05085e56",
972 => x"7c762e84",
973 => x"bd388416",
974 => x"0870fe06",
975 => x"17841108",
976 => x"81065155",
977 => x"5573828b",
978 => x"3874fc06",
979 => x"597c762e",
980 => x"84dd3877",
981 => x"195f7e7b",
982 => x"2581fd38",
983 => x"79810654",
984 => x"7382bf38",
985 => x"76770831",
986 => x"841108fc",
987 => x"06565a75",
988 => x"802e9138",
989 => x"7c762e84",
990 => x"ea387419",
991 => x"1859787b",
992 => x"25848938",
993 => x"79802e82",
994 => x"99387715",
995 => x"567a7624",
996 => x"8290388c",
997 => x"1a08881b",
998 => x"08718c12",
999 => x"0c88120c",
1000 => x"55797659",
1001 => x"57881761",
1002 => x"fc055759",
1003 => x"75a42685",
1004 => x"ef387b79",
1005 => x"55559376",
1006 => x"2780c938",
1007 => x"7b708405",
1008 => x"5d087c56",
1009 => x"790c7470",
1010 => x"84055608",
1011 => x"8c180c90",
1012 => x"17549b76",
1013 => x"27ae3874",
1014 => x"70840556",
1015 => x"08740c74",
1016 => x"70840556",
1017 => x"0894180c",
1018 => x"981754a3",
1019 => x"76279538",
1020 => x"74708405",
1021 => x"5608740c",
1022 => x"74708405",
1023 => x"56089c18",
1024 => x"0ca01754",
1025 => x"74708405",
1026 => x"56087470",
1027 => x"8405560c",
1028 => x"74708405",
1029 => x"56087470",
1030 => x"8405560c",
1031 => x"7408740c",
1032 => x"777b3156",
1033 => x"758f2680",
1034 => x"c9388417",
1035 => x"08810678",
1036 => x"0784180c",
1037 => x"77178411",
1038 => x"08810784",
1039 => x"120c5461",
1040 => x"51a2e03f",
1041 => x"88175473",
1042 => x"b00c933d",
1043 => x"0d04905b",
1044 => x"fdba3978",
1045 => x"56fe8539",
1046 => x"8c160888",
1047 => x"1708718c",
1048 => x"120c8812",
1049 => x"0c557e70",
1050 => x"7c315758",
1051 => x"8f7627ff",
1052 => x"b9387a17",
1053 => x"84180881",
1054 => x"067c0784",
1055 => x"190c7681",
1056 => x"0784120c",
1057 => x"76118411",
1058 => x"08810784",
1059 => x"120c5588",
1060 => x"05526151",
1061 => x"8cf63f61",
1062 => x"51a2883f",
1063 => x"881754ff",
1064 => x"a6397d52",
1065 => x"615194f5",
1066 => x"3fb00859",
1067 => x"b008802e",
1068 => x"81a338b0",
1069 => x"08f80560",
1070 => x"840508fe",
1071 => x"06610555",
1072 => x"5776742e",
1073 => x"83e638fc",
1074 => x"185675a4",
1075 => x"2681aa38",
1076 => x"7bb00855",
1077 => x"55937627",
1078 => x"80d83874",
1079 => x"70840556",
1080 => x"08b00870",
1081 => x"8405b00c",
1082 => x"0cb00875",
1083 => x"70840557",
1084 => x"08717084",
1085 => x"05530c54",
1086 => x"9b7627b6",
1087 => x"38747084",
1088 => x"05560874",
1089 => x"70840556",
1090 => x"0c747084",
1091 => x"05560874",
1092 => x"70840556",
1093 => x"0ca37627",
1094 => x"99387470",
1095 => x"84055608",
1096 => x"74708405",
1097 => x"560c7470",
1098 => x"84055608",
1099 => x"74708405",
1100 => x"560c7470",
1101 => x"84055608",
1102 => x"74708405",
1103 => x"560c7470",
1104 => x"84055608",
1105 => x"74708405",
1106 => x"560c7408",
1107 => x"740c7b52",
1108 => x"61518bb8",
1109 => x"3f6151a0",
1110 => x"ca3f7854",
1111 => x"73b00c93",
1112 => x"3d0d047d",
1113 => x"52615193",
1114 => x"b43fb008",
1115 => x"b00c933d",
1116 => x"0d048416",
1117 => x"0855fbd1",
1118 => x"3975537b",
1119 => x"52b00851",
1120 => x"efc63f7b",
1121 => x"5261518b",
1122 => x"833fca39",
1123 => x"8c160888",
1124 => x"1708718c",
1125 => x"120c8812",
1126 => x"0c558c1a",
1127 => x"08881b08",
1128 => x"718c120c",
1129 => x"88120c55",
1130 => x"79795957",
1131 => x"fbf73977",
1132 => x"19901c55",
1133 => x"55737524",
1134 => x"fba2387a",
1135 => x"177080d8",
1136 => x"c00b8805",
1137 => x"0c757c31",
1138 => x"81078412",
1139 => x"0c5d8417",
1140 => x"0881067b",
1141 => x"0784180c",
1142 => x"61519fc7",
1143 => x"3f881754",
1144 => x"fce53974",
1145 => x"1918901c",
1146 => x"555d737d",
1147 => x"24fb9538",
1148 => x"8c1a0888",
1149 => x"1b08718c",
1150 => x"120c8812",
1151 => x"0c55881a",
1152 => x"61fc0557",
1153 => x"5975a426",
1154 => x"81ae387b",
1155 => x"79555593",
1156 => x"762780c9",
1157 => x"387b7084",
1158 => x"055d087c",
1159 => x"56790c74",
1160 => x"70840556",
1161 => x"088c1b0c",
1162 => x"901a549b",
1163 => x"7627ae38",
1164 => x"74708405",
1165 => x"5608740c",
1166 => x"74708405",
1167 => x"5608941b",
1168 => x"0c981a54",
1169 => x"a3762795",
1170 => x"38747084",
1171 => x"05560874",
1172 => x"0c747084",
1173 => x"0556089c",
1174 => x"1b0ca01a",
1175 => x"54747084",
1176 => x"05560874",
1177 => x"70840556",
1178 => x"0c747084",
1179 => x"05560874",
1180 => x"70840556",
1181 => x"0c740874",
1182 => x"0c7a1a70",
1183 => x"80d8c00b",
1184 => x"88050c7d",
1185 => x"7c318107",
1186 => x"84120c54",
1187 => x"841a0881",
1188 => x"067b0784",
1189 => x"1b0c6151",
1190 => x"9e893f78",
1191 => x"54fdbd39",
1192 => x"75537b52",
1193 => x"7851eda0",
1194 => x"3ffaf539",
1195 => x"841708fc",
1196 => x"06186058",
1197 => x"58fae939",
1198 => x"75537b52",
1199 => x"7851ed88",
1200 => x"3f7a1a70",
1201 => x"80d8c00b",
1202 => x"88050c7d",
1203 => x"7c318107",
1204 => x"84120c54",
1205 => x"841a0881",
1206 => x"067b0784",
1207 => x"1b0cffb6",
1208 => x"39fa3d0d",
1209 => x"7880d184",
1210 => x"085455b8",
1211 => x"1308802e",
1212 => x"81b5388c",
1213 => x"15227083",
1214 => x"ffff0670",
1215 => x"832a8132",
1216 => x"70810651",
1217 => x"55555672",
1218 => x"802e80dc",
1219 => x"3873842a",
1220 => x"81328106",
1221 => x"57ff5376",
1222 => x"80f63873",
1223 => x"822a7081",
1224 => x"06515372",
1225 => x"802eb938",
1226 => x"b0150854",
1227 => x"73802e9c",
1228 => x"3880c015",
1229 => x"5373732e",
1230 => x"8f387352",
1231 => x"80d18408",
1232 => x"5187c93f",
1233 => x"8c152256",
1234 => x"76b0160c",
1235 => x"75db0653",
1236 => x"728c1623",
1237 => x"800b8416",
1238 => x"0c901508",
1239 => x"750c7256",
1240 => x"75880753",
1241 => x"728c1623",
1242 => x"90150880",
1243 => x"2e80c038",
1244 => x"8c152270",
1245 => x"81065553",
1246 => x"739d3872",
1247 => x"812a7081",
1248 => x"06515372",
1249 => x"85389415",
1250 => x"08547388",
1251 => x"160c8053",
1252 => x"72b00c88",
1253 => x"3d0d0480",
1254 => x"0b88160c",
1255 => x"94150830",
1256 => x"98160c80",
1257 => x"53ea3972",
1258 => x"5182fb3f",
1259 => x"fec53974",
1260 => x"518ce83f",
1261 => x"8c152270",
1262 => x"81065553",
1263 => x"73802eff",
1264 => x"ba38d439",
1265 => x"f83d0d7a",
1266 => x"5877802e",
1267 => x"81993880",
1268 => x"d1840854",
1269 => x"b8140880",
1270 => x"2e80ed38",
1271 => x"8c182270",
1272 => x"902b7090",
1273 => x"2c70832a",
1274 => x"81328106",
1275 => x"5c515754",
1276 => x"7880cd38",
1277 => x"90180857",
1278 => x"76802e80",
1279 => x"c3387708",
1280 => x"77317779",
1281 => x"0c768306",
1282 => x"7a585555",
1283 => x"73853894",
1284 => x"18085675",
1285 => x"88190c80",
1286 => x"7525a538",
1287 => x"74537652",
1288 => x"9c180851",
1289 => x"a4180854",
1290 => x"732d800b",
1291 => x"b0082580",
1292 => x"c938b008",
1293 => x"1775b008",
1294 => x"31565774",
1295 => x"8024dd38",
1296 => x"800bb00c",
1297 => x"8a3d0d04",
1298 => x"735181da",
1299 => x"3f8c1822",
1300 => x"70902b70",
1301 => x"902c7083",
1302 => x"2a813281",
1303 => x"065c5157",
1304 => x"5478dd38",
1305 => x"ff8e39a7",
1306 => x"c45280d1",
1307 => x"84085189",
1308 => x"f13fb008",
1309 => x"b00c8a3d",
1310 => x"0d048c18",
1311 => x"2280c007",
1312 => x"54738c19",
1313 => x"23ff0bb0",
1314 => x"0c8a3d0d",
1315 => x"04803d0d",
1316 => x"72518071",
1317 => x"0c800b84",
1318 => x"120c800b",
1319 => x"88120c02",
1320 => x"8e05228c",
1321 => x"12230292",
1322 => x"05228e12",
1323 => x"23800b90",
1324 => x"120c800b",
1325 => x"94120c80",
1326 => x"0b98120c",
1327 => x"709c120c",
1328 => x"80c3d80b",
1329 => x"a0120c80",
1330 => x"c4a40ba4",
1331 => x"120c80c5",
1332 => x"a00ba812",
1333 => x"0c80c5f1",
1334 => x"0bac120c",
1335 => x"823d0d04",
1336 => x"fa3d0d79",
1337 => x"7080dc29",
1338 => x"8c11547a",
1339 => x"5356578c",
1340 => x"ac3fb008",
1341 => x"b0085556",
1342 => x"b008802e",
1343 => x"a238b008",
1344 => x"8c055480",
1345 => x"0bb0080c",
1346 => x"76b00884",
1347 => x"050c73b0",
1348 => x"0888050c",
1349 => x"74538052",
1350 => x"735197f7",
1351 => x"3f755473",
1352 => x"b00c883d",
1353 => x"0d04fc3d",
1354 => x"0d76acb9",
1355 => x"0bbc120c",
1356 => x"55810bb8",
1357 => x"160c800b",
1358 => x"84dc160c",
1359 => x"830b84e0",
1360 => x"160c84e8",
1361 => x"1584e416",
1362 => x"0c745480",
1363 => x"53845284",
1364 => x"150851fe",
1365 => x"b83f7454",
1366 => x"81538952",
1367 => x"88150851",
1368 => x"feab3f74",
1369 => x"5482538a",
1370 => x"528c1508",
1371 => x"51fe9e3f",
1372 => x"863d0d04",
1373 => x"f93d0d79",
1374 => x"80d18408",
1375 => x"5457b813",
1376 => x"08802e80",
1377 => x"c83884dc",
1378 => x"13568816",
1379 => x"08841708",
1380 => x"ff055555",
1381 => x"8074249f",
1382 => x"388c1522",
1383 => x"70902b70",
1384 => x"902c5154",
1385 => x"5872802e",
1386 => x"80ca3880",
1387 => x"dc15ff15",
1388 => x"55557380",
1389 => x"25e33875",
1390 => x"08537280",
1391 => x"2e9f3872",
1392 => x"56881608",
1393 => x"841708ff",
1394 => x"055555c8",
1395 => x"397251fe",
1396 => x"d53f80d1",
1397 => x"840884dc",
1398 => x"0556ffae",
1399 => x"39845276",
1400 => x"51fdfd3f",
1401 => x"b008760c",
1402 => x"b008802e",
1403 => x"80c038b0",
1404 => x"0856ce39",
1405 => x"810b8c16",
1406 => x"2372750c",
1407 => x"7288160c",
1408 => x"7284160c",
1409 => x"7290160c",
1410 => x"7294160c",
1411 => x"7298160c",
1412 => x"ff0b8e16",
1413 => x"2372b016",
1414 => x"0c72b416",
1415 => x"0c7280c4",
1416 => x"160c7280",
1417 => x"c8160c74",
1418 => x"b00c893d",
1419 => x"0d048c77",
1420 => x"0c800bb0",
1421 => x"0c893d0d",
1422 => x"04ff3d0d",
1423 => x"a7c45273",
1424 => x"51869f3f",
1425 => x"833d0d04",
1426 => x"803d0d80",
1427 => x"d1840851",
1428 => x"e83f823d",
1429 => x"0d04fb3d",
1430 => x"0d777052",
1431 => x"5696c33f",
1432 => x"80d8c00b",
1433 => x"88050884",
1434 => x"1108fc06",
1435 => x"707b319f",
1436 => x"ef05e080",
1437 => x"06e08005",
1438 => x"565653a0",
1439 => x"80742494",
1440 => x"38805275",
1441 => x"51969d3f",
1442 => x"80d8c808",
1443 => x"155372b0",
1444 => x"082e8f38",
1445 => x"7551968b",
1446 => x"3f805372",
1447 => x"b00c873d",
1448 => x"0d047330",
1449 => x"52755195",
1450 => x"fb3fb008",
1451 => x"ff2ea838",
1452 => x"80d8c00b",
1453 => x"88050875",
1454 => x"75318107",
1455 => x"84120c53",
1456 => x"80d88408",
1457 => x"743180d8",
1458 => x"840c7551",
1459 => x"95d53f81",
1460 => x"0bb00c87",
1461 => x"3d0d0480",
1462 => x"52755195",
1463 => x"c73f80d8",
1464 => x"c00b8805",
1465 => x"08b00871",
1466 => x"3156538f",
1467 => x"7525ffa4",
1468 => x"38b00880",
1469 => x"d8b40831",
1470 => x"80d8840c",
1471 => x"74810784",
1472 => x"140c7551",
1473 => x"959d3f80",
1474 => x"53ff9039",
1475 => x"f63d0d7c",
1476 => x"7e545b72",
1477 => x"802e8283",
1478 => x"387a5195",
1479 => x"853ff813",
1480 => x"84110870",
1481 => x"fe067013",
1482 => x"841108fc",
1483 => x"065d5859",
1484 => x"545880d8",
1485 => x"c808752e",
1486 => x"82de3878",
1487 => x"84160c80",
1488 => x"73810654",
1489 => x"5a727a2e",
1490 => x"81d53878",
1491 => x"15841108",
1492 => x"81065153",
1493 => x"72a03878",
1494 => x"17577981",
1495 => x"e6388815",
1496 => x"08537280",
1497 => x"d8c82e82",
1498 => x"f9388c15",
1499 => x"08708c15",
1500 => x"0c738812",
1501 => x"0c567681",
1502 => x"0784190c",
1503 => x"76187771",
1504 => x"0c537981",
1505 => x"913883ff",
1506 => x"772781c8",
1507 => x"3876892a",
1508 => x"77832a56",
1509 => x"5372802e",
1510 => x"bf387686",
1511 => x"2ab80555",
1512 => x"847327b4",
1513 => x"3880db13",
1514 => x"55947327",
1515 => x"ab38768c",
1516 => x"2a80ee05",
1517 => x"5580d473",
1518 => x"279e3876",
1519 => x"8f2a80f7",
1520 => x"055582d4",
1521 => x"73279138",
1522 => x"76922a80",
1523 => x"fc05558a",
1524 => x"d4732784",
1525 => x"3880fe55",
1526 => x"74101010",
1527 => x"80d8c005",
1528 => x"88110855",
1529 => x"5673762e",
1530 => x"82b33884",
1531 => x"1408fc06",
1532 => x"53767327",
1533 => x"8d388814",
1534 => x"08547376",
1535 => x"2e098106",
1536 => x"ea388c14",
1537 => x"08708c1a",
1538 => x"0c74881a",
1539 => x"0c788812",
1540 => x"0c56778c",
1541 => x"150c7a51",
1542 => x"93893f8c",
1543 => x"3d0d0477",
1544 => x"08787131",
1545 => x"59770588",
1546 => x"19085457",
1547 => x"7280d8c8",
1548 => x"2e80e038",
1549 => x"8c180870",
1550 => x"8c150c73",
1551 => x"88120c56",
1552 => x"fe893988",
1553 => x"15088c16",
1554 => x"08708c13",
1555 => x"0c578817",
1556 => x"0cfea339",
1557 => x"76832a70",
1558 => x"54558075",
1559 => x"24819838",
1560 => x"72822c81",
1561 => x"712b80d8",
1562 => x"c4080780",
1563 => x"d8c00b84",
1564 => x"050c5374",
1565 => x"10101080",
1566 => x"d8c00588",
1567 => x"11085556",
1568 => x"758c190c",
1569 => x"7388190c",
1570 => x"7788170c",
1571 => x"778c150c",
1572 => x"ff843981",
1573 => x"5afdb439",
1574 => x"78177381",
1575 => x"06545772",
1576 => x"98387708",
1577 => x"78713159",
1578 => x"77058c19",
1579 => x"08881a08",
1580 => x"718c120c",
1581 => x"88120c57",
1582 => x"57768107",
1583 => x"84190c77",
1584 => x"80d8c00b",
1585 => x"88050c80",
1586 => x"d8bc0877",
1587 => x"26fec738",
1588 => x"80d8b808",
1589 => x"527a51fa",
1590 => x"fd3f7a51",
1591 => x"91c53ffe",
1592 => x"ba398178",
1593 => x"8c150c78",
1594 => x"88150c73",
1595 => x"8c1a0c73",
1596 => x"881a0c5a",
1597 => x"fd803983",
1598 => x"1570822c",
1599 => x"81712b80",
1600 => x"d8c40807",
1601 => x"80d8c00b",
1602 => x"84050c51",
1603 => x"53741010",
1604 => x"1080d8c0",
1605 => x"05881108",
1606 => x"5556fee4",
1607 => x"39745380",
1608 => x"7524a738",
1609 => x"72822c81",
1610 => x"712b80d8",
1611 => x"c4080780",
1612 => x"d8c00b84",
1613 => x"050c5375",
1614 => x"8c190c73",
1615 => x"88190c77",
1616 => x"88170c77",
1617 => x"8c150cfd",
1618 => x"cd398315",
1619 => x"70822c81",
1620 => x"712b80d8",
1621 => x"c4080780",
1622 => x"d8c00b84",
1623 => x"050c5153",
1624 => x"d639f93d",
1625 => x"0d797b58",
1626 => x"53800b80",
1627 => x"d1840853",
1628 => x"5672722e",
1629 => x"80c03884",
1630 => x"dc135574",
1631 => x"762eb738",
1632 => x"88150884",
1633 => x"1608ff05",
1634 => x"54548073",
1635 => x"249d388c",
1636 => x"14227090",
1637 => x"2b70902c",
1638 => x"51535871",
1639 => x"80d83880",
1640 => x"dc14ff14",
1641 => x"54547280",
1642 => x"25e53874",
1643 => x"085574d0",
1644 => x"3880d184",
1645 => x"085284dc",
1646 => x"12557480",
1647 => x"2eb13888",
1648 => x"15088416",
1649 => x"08ff0554",
1650 => x"54807324",
1651 => x"9c388c14",
1652 => x"2270902b",
1653 => x"70902c51",
1654 => x"535871ad",
1655 => x"3880dc14",
1656 => x"ff145454",
1657 => x"728025e6",
1658 => x"38740855",
1659 => x"74d13875",
1660 => x"b00c893d",
1661 => x"0d047351",
1662 => x"762d75b0",
1663 => x"080780dc",
1664 => x"15ff1555",
1665 => x"5556ff9e",
1666 => x"39735176",
1667 => x"2d75b008",
1668 => x"0780dc15",
1669 => x"ff155555",
1670 => x"56ca39ea",
1671 => x"3d0d688c",
1672 => x"11227081",
1673 => x"2a810657",
1674 => x"58567480",
1675 => x"e4388e16",
1676 => x"2270902b",
1677 => x"70902c51",
1678 => x"55588074",
1679 => x"24b13898",
1680 => x"3dc40553",
1681 => x"735280d1",
1682 => x"84085192",
1683 => x"ac3f800b",
1684 => x"b0082497",
1685 => x"387983e0",
1686 => x"80065473",
1687 => x"80c0802e",
1688 => x"818f3873",
1689 => x"8280802e",
1690 => x"8191388c",
1691 => x"16225776",
1692 => x"90800754",
1693 => x"738c1723",
1694 => x"88805280",
1695 => x"d1840851",
1696 => x"819b3fb0",
1697 => x"089d388c",
1698 => x"16228207",
1699 => x"54738c17",
1700 => x"2380c316",
1701 => x"70770c90",
1702 => x"170c810b",
1703 => x"94170c98",
1704 => x"3d0d0480",
1705 => x"d18408ac",
1706 => x"b90bbc12",
1707 => x"0c548c16",
1708 => x"22818007",
1709 => x"54738c17",
1710 => x"23b00876",
1711 => x"0cb00890",
1712 => x"170c8880",
1713 => x"0b94170c",
1714 => x"74802ed3",
1715 => x"388e1622",
1716 => x"70902b70",
1717 => x"902c5355",
1718 => x"5898ae3f",
1719 => x"b008802e",
1720 => x"ffbd388c",
1721 => x"16228107",
1722 => x"54738c17",
1723 => x"23983d0d",
1724 => x"04810b8c",
1725 => x"17225855",
1726 => x"fef539a8",
1727 => x"160880c5",
1728 => x"a02e0981",
1729 => x"06fee438",
1730 => x"8c162288",
1731 => x"80075473",
1732 => x"8c172388",
1733 => x"800b80cc",
1734 => x"170cfedc",
1735 => x"39f33d0d",
1736 => x"7f618b11",
1737 => x"70f8065c",
1738 => x"55555e72",
1739 => x"96268338",
1740 => x"90598079",
1741 => x"24747a26",
1742 => x"07538054",
1743 => x"72742e09",
1744 => x"810680cb",
1745 => x"387d518c",
1746 => x"d93f7883",
1747 => x"f72680c6",
1748 => x"3878832a",
1749 => x"70101010",
1750 => x"80d8c005",
1751 => x"8c110859",
1752 => x"595a7678",
1753 => x"2e83b038",
1754 => x"841708fc",
1755 => x"06568c17",
1756 => x"08881808",
1757 => x"718c120c",
1758 => x"88120c58",
1759 => x"75178411",
1760 => x"08810784",
1761 => x"120c537d",
1762 => x"518c983f",
1763 => x"88175473",
1764 => x"b00c8f3d",
1765 => x"0d047889",
1766 => x"2a79832a",
1767 => x"5b537280",
1768 => x"2ebf3878",
1769 => x"862ab805",
1770 => x"5a847327",
1771 => x"b43880db",
1772 => x"135a9473",
1773 => x"27ab3878",
1774 => x"8c2a80ee",
1775 => x"055a80d4",
1776 => x"73279e38",
1777 => x"788f2a80",
1778 => x"f7055a82",
1779 => x"d4732791",
1780 => x"3878922a",
1781 => x"80fc055a",
1782 => x"8ad47327",
1783 => x"843880fe",
1784 => x"5a791010",
1785 => x"1080d8c0",
1786 => x"058c1108",
1787 => x"58557675",
1788 => x"2ea33884",
1789 => x"1708fc06",
1790 => x"707a3155",
1791 => x"56738f24",
1792 => x"88d53873",
1793 => x"8025fee6",
1794 => x"388c1708",
1795 => x"5776752e",
1796 => x"098106df",
1797 => x"38811a5a",
1798 => x"80d8d008",
1799 => x"577680d8",
1800 => x"c82e82c0",
1801 => x"38841708",
1802 => x"fc06707a",
1803 => x"31555673",
1804 => x"8f2481f9",
1805 => x"3880d8c8",
1806 => x"0b80d8d4",
1807 => x"0c80d8c8",
1808 => x"0b80d8d0",
1809 => x"0c738025",
1810 => x"feb23883",
1811 => x"ff762783",
1812 => x"df387589",
1813 => x"2a76832a",
1814 => x"55537280",
1815 => x"2ebf3875",
1816 => x"862ab805",
1817 => x"54847327",
1818 => x"b43880db",
1819 => x"13549473",
1820 => x"27ab3875",
1821 => x"8c2a80ee",
1822 => x"055480d4",
1823 => x"73279e38",
1824 => x"758f2a80",
1825 => x"f7055482",
1826 => x"d4732791",
1827 => x"3875922a",
1828 => x"80fc0554",
1829 => x"8ad47327",
1830 => x"843880fe",
1831 => x"54731010",
1832 => x"1080d8c0",
1833 => x"05881108",
1834 => x"56587478",
1835 => x"2e86cf38",
1836 => x"841508fc",
1837 => x"06537573",
1838 => x"278d3888",
1839 => x"15085574",
1840 => x"782e0981",
1841 => x"06ea388c",
1842 => x"150880d8",
1843 => x"c00b8405",
1844 => x"08718c1a",
1845 => x"0c76881a",
1846 => x"0c788813",
1847 => x"0c788c18",
1848 => x"0c5d5879",
1849 => x"53807a24",
1850 => x"83e63872",
1851 => x"822c8171",
1852 => x"2b5c537a",
1853 => x"7c268198",
1854 => x"387b7b06",
1855 => x"537282f1",
1856 => x"3879fc06",
1857 => x"84055a7a",
1858 => x"10707d06",
1859 => x"545b7282",
1860 => x"e038841a",
1861 => x"5af13988",
1862 => x"178c1108",
1863 => x"58587678",
1864 => x"2e098106",
1865 => x"fcc23882",
1866 => x"1a5afdec",
1867 => x"39781779",
1868 => x"81078419",
1869 => x"0c7080d8",
1870 => x"d40c7080",
1871 => x"d8d00c80",
1872 => x"d8c80b8c",
1873 => x"120c8c11",
1874 => x"0888120c",
1875 => x"74810784",
1876 => x"120c7411",
1877 => x"75710c51",
1878 => x"537d5188",
1879 => x"c63f8817",
1880 => x"54fcac39",
1881 => x"80d8c00b",
1882 => x"8405087a",
1883 => x"545c7980",
1884 => x"25fef838",
1885 => x"82da397a",
1886 => x"097c0670",
1887 => x"80d8c00b",
1888 => x"84050c5c",
1889 => x"7a105b7a",
1890 => x"7c268538",
1891 => x"7a85b838",
1892 => x"80d8c00b",
1893 => x"88050870",
1894 => x"841208fc",
1895 => x"06707c31",
1896 => x"7c72268f",
1897 => x"72250757",
1898 => x"575c5d55",
1899 => x"72802e80",
1900 => x"db38797a",
1901 => x"1680d8b8",
1902 => x"081b9011",
1903 => x"5a55575b",
1904 => x"80d8b408",
1905 => x"ff2e8838",
1906 => x"a08f13e0",
1907 => x"80065776",
1908 => x"527d5187",
1909 => x"cf3fb008",
1910 => x"54b008ff",
1911 => x"2e9038b0",
1912 => x"08762782",
1913 => x"99387480",
1914 => x"d8c02e82",
1915 => x"913880d8",
1916 => x"c00b8805",
1917 => x"08558415",
1918 => x"08fc0670",
1919 => x"7a317a72",
1920 => x"268f7225",
1921 => x"07525553",
1922 => x"7283e638",
1923 => x"74798107",
1924 => x"84170c79",
1925 => x"167080d8",
1926 => x"c00b8805",
1927 => x"0c758107",
1928 => x"84120c54",
1929 => x"7e525786",
1930 => x"fa3f8817",
1931 => x"54fae039",
1932 => x"75832a70",
1933 => x"54548074",
1934 => x"24819b38",
1935 => x"72822c81",
1936 => x"712b80d8",
1937 => x"c4080770",
1938 => x"80d8c00b",
1939 => x"84050c75",
1940 => x"10101080",
1941 => x"d8c00588",
1942 => x"1108585a",
1943 => x"5d53778c",
1944 => x"180c7488",
1945 => x"180c7688",
1946 => x"190c768c",
1947 => x"160cfcf3",
1948 => x"39797a10",
1949 => x"101080d8",
1950 => x"c0057057",
1951 => x"595d8c15",
1952 => x"08577675",
1953 => x"2ea33884",
1954 => x"1708fc06",
1955 => x"707a3155",
1956 => x"56738f24",
1957 => x"83ca3873",
1958 => x"80258481",
1959 => x"388c1708",
1960 => x"5776752e",
1961 => x"098106df",
1962 => x"38881581",
1963 => x"1b708306",
1964 => x"555b5572",
1965 => x"c9387c83",
1966 => x"06537280",
1967 => x"2efdb838",
1968 => x"ff1df819",
1969 => x"595d8818",
1970 => x"08782eea",
1971 => x"38fdb539",
1972 => x"831a53fc",
1973 => x"96398314",
1974 => x"70822c81",
1975 => x"712b80d8",
1976 => x"c4080770",
1977 => x"80d8c00b",
1978 => x"84050c76",
1979 => x"10101080",
1980 => x"d8c00588",
1981 => x"1108595b",
1982 => x"5e5153fe",
1983 => x"e13980d8",
1984 => x"84081758",
1985 => x"b008762e",
1986 => x"818d3880",
1987 => x"d8b408ff",
1988 => x"2e83ec38",
1989 => x"73763118",
1990 => x"80d8840c",
1991 => x"73870670",
1992 => x"57537280",
1993 => x"2e883888",
1994 => x"73317015",
1995 => x"55567614",
1996 => x"9fff06a0",
1997 => x"80713117",
1998 => x"70547f53",
1999 => x"575384e4",
2000 => x"3fb00853",
2001 => x"b008ff2e",
2002 => x"81a03880",
2003 => x"d8840816",
2004 => x"7080d884",
2005 => x"0c747580",
2006 => x"d8c00b88",
2007 => x"050c7476",
2008 => x"31187081",
2009 => x"07515556",
2010 => x"587b80d8",
2011 => x"c02e839c",
2012 => x"38798f26",
2013 => x"82cb3881",
2014 => x"0b84150c",
2015 => x"841508fc",
2016 => x"06707a31",
2017 => x"7a72268f",
2018 => x"72250752",
2019 => x"55537280",
2020 => x"2efcf938",
2021 => x"80db39b0",
2022 => x"089fff06",
2023 => x"5372feeb",
2024 => x"387780d8",
2025 => x"840c80d8",
2026 => x"c00b8805",
2027 => x"087b1881",
2028 => x"0784120c",
2029 => x"5580d8b0",
2030 => x"08782786",
2031 => x"387780d8",
2032 => x"b00c80d8",
2033 => x"ac087827",
2034 => x"fcac3877",
2035 => x"80d8ac0c",
2036 => x"841508fc",
2037 => x"06707a31",
2038 => x"7a72268f",
2039 => x"72250752",
2040 => x"55537280",
2041 => x"2efca538",
2042 => x"88398074",
2043 => x"5456fedb",
2044 => x"397d5183",
2045 => x"ae3f800b",
2046 => x"b00c8f3d",
2047 => x"0d047353",
2048 => x"807424a9",
2049 => x"3872822c",
2050 => x"81712b80",
2051 => x"d8c40807",
2052 => x"7080d8c0",
2053 => x"0b84050c",
2054 => x"5d53778c",
2055 => x"180c7488",
2056 => x"180c7688",
2057 => x"190c768c",
2058 => x"160cf9b7",
2059 => x"39831470",
2060 => x"822c8171",
2061 => x"2b80d8c4",
2062 => x"08077080",
2063 => x"d8c00b84",
2064 => x"050c5e51",
2065 => x"53d4397b",
2066 => x"7b065372",
2067 => x"fca33884",
2068 => x"1a7b105c",
2069 => x"5af139ff",
2070 => x"1a811151",
2071 => x"5af7b939",
2072 => x"78177981",
2073 => x"0784190c",
2074 => x"8c180888",
2075 => x"1908718c",
2076 => x"120c8812",
2077 => x"0c597080",
2078 => x"d8d40c70",
2079 => x"80d8d00c",
2080 => x"80d8c80b",
2081 => x"8c120c8c",
2082 => x"11088812",
2083 => x"0c748107",
2084 => x"84120c74",
2085 => x"1175710c",
2086 => x"5153f9bd",
2087 => x"39751784",
2088 => x"11088107",
2089 => x"84120c53",
2090 => x"8c170888",
2091 => x"1808718c",
2092 => x"120c8812",
2093 => x"0c587d51",
2094 => x"81e93f88",
2095 => x"1754f5cf",
2096 => x"39728415",
2097 => x"0cf41af8",
2098 => x"0670841e",
2099 => x"08810607",
2100 => x"841e0c70",
2101 => x"1d545b85",
2102 => x"0b84140c",
2103 => x"850b8814",
2104 => x"0c8f7b27",
2105 => x"fdcf3888",
2106 => x"1c527d51",
2107 => x"ec9e3f80",
2108 => x"d8c00b88",
2109 => x"050880d8",
2110 => x"84085955",
2111 => x"fdb73977",
2112 => x"80d8840c",
2113 => x"7380d8b4",
2114 => x"0cfc9139",
2115 => x"7284150c",
2116 => x"fda339fc",
2117 => x"3d0d7679",
2118 => x"71028c05",
2119 => x"9f053357",
2120 => x"55535583",
2121 => x"72278a38",
2122 => x"74830651",
2123 => x"70802ea2",
2124 => x"38ff1252",
2125 => x"71ff2e93",
2126 => x"38737370",
2127 => x"81055534",
2128 => x"ff125271",
2129 => x"ff2e0981",
2130 => x"06ef3874",
2131 => x"b00c863d",
2132 => x"0d047474",
2133 => x"882b7507",
2134 => x"7071902b",
2135 => x"07515451",
2136 => x"8f7227a5",
2137 => x"38727170",
2138 => x"8405530c",
2139 => x"72717084",
2140 => x"05530c72",
2141 => x"71708405",
2142 => x"530c7271",
2143 => x"70840553",
2144 => x"0cf01252",
2145 => x"718f26dd",
2146 => x"38837227",
2147 => x"90387271",
2148 => x"70840553",
2149 => x"0cfc1252",
2150 => x"718326f2",
2151 => x"387053ff",
2152 => x"90390404",
2153 => x"fd3d0d80",
2154 => x"0b80e0fc",
2155 => x"0c765184",
2156 => x"ee3fb008",
2157 => x"53b008ff",
2158 => x"2e883872",
2159 => x"b00c853d",
2160 => x"0d0480e0",
2161 => x"fc085473",
2162 => x"802ef038",
2163 => x"7574710c",
2164 => x"5272b00c",
2165 => x"853d0d04",
2166 => x"f93d0d79",
2167 => x"7c557b54",
2168 => x"8e112270",
2169 => x"902b7090",
2170 => x"2c555780",
2171 => x"d1840853",
2172 => x"585683f3",
2173 => x"3fb00857",
2174 => x"800bb008",
2175 => x"24933880",
2176 => x"d01608b0",
2177 => x"080580d0",
2178 => x"170c76b0",
2179 => x"0c893d0d",
2180 => x"048c1622",
2181 => x"83dfff06",
2182 => x"55748c17",
2183 => x"2376b00c",
2184 => x"893d0d04",
2185 => x"fa3d0d78",
2186 => x"8c112270",
2187 => x"882a7081",
2188 => x"06515758",
2189 => x"5674a938",
2190 => x"8c162283",
2191 => x"dfff0655",
2192 => x"748c1723",
2193 => x"7a547953",
2194 => x"8e162270",
2195 => x"902b7090",
2196 => x"2c545680",
2197 => x"d1840852",
2198 => x"5681b23f",
2199 => x"883d0d04",
2200 => x"82548053",
2201 => x"8e162270",
2202 => x"902b7090",
2203 => x"2c545680",
2204 => x"d1840852",
2205 => x"5782b83f",
2206 => x"8c162283",
2207 => x"dfff0655",
2208 => x"748c1723",
2209 => x"7a547953",
2210 => x"8e162270",
2211 => x"902b7090",
2212 => x"2c545680",
2213 => x"d1840852",
2214 => x"5680f23f",
2215 => x"883d0d04",
2216 => x"f93d0d79",
2217 => x"7c557b54",
2218 => x"8e112270",
2219 => x"902b7090",
2220 => x"2c555780",
2221 => x"d1840853",
2222 => x"585681f3",
2223 => x"3fb00857",
2224 => x"b008ff2e",
2225 => x"99388c16",
2226 => x"22a08007",
2227 => x"55748c17",
2228 => x"23b00880",
2229 => x"d0170c76",
2230 => x"b00c893d",
2231 => x"0d048c16",
2232 => x"2283dfff",
2233 => x"0655748c",
2234 => x"172376b0",
2235 => x"0c893d0d",
2236 => x"04fe3d0d",
2237 => x"748e1122",
2238 => x"70902b70",
2239 => x"902c5551",
2240 => x"515380d1",
2241 => x"840851bd",
2242 => x"3f843d0d",
2243 => x"04fb3d0d",
2244 => x"800b80e0",
2245 => x"fc0c7a53",
2246 => x"79527851",
2247 => x"82fb3fb0",
2248 => x"0855b008",
2249 => x"ff2e8838",
2250 => x"74b00c87",
2251 => x"3d0d0480",
2252 => x"e0fc0856",
2253 => x"75802ef0",
2254 => x"38777671",
2255 => x"0c5474b0",
2256 => x"0c873d0d",
2257 => x"04fd3d0d",
2258 => x"800b80e0",
2259 => x"fc0c7651",
2260 => x"84d03fb0",
2261 => x"0853b008",
2262 => x"ff2e8838",
2263 => x"72b00c85",
2264 => x"3d0d0480",
2265 => x"e0fc0854",
2266 => x"73802ef0",
2267 => x"38757471",
2268 => x"0c5272b0",
2269 => x"0c853d0d",
2270 => x"04fc3d0d",
2271 => x"800b80e0",
2272 => x"fc0c7852",
2273 => x"775186b8",
2274 => x"3fb00854",
2275 => x"b008ff2e",
2276 => x"883873b0",
2277 => x"0c863d0d",
2278 => x"0480e0fc",
2279 => x"08557480",
2280 => x"2ef03876",
2281 => x"75710c53",
2282 => x"73b00c86",
2283 => x"3d0d04fb",
2284 => x"3d0d800b",
2285 => x"80e0fc0c",
2286 => x"7a537952",
2287 => x"78518494",
2288 => x"3fb00855",
2289 => x"b008ff2e",
2290 => x"883874b0",
2291 => x"0c873d0d",
2292 => x"0480e0fc",
2293 => x"08567580",
2294 => x"2ef03877",
2295 => x"76710c54",
2296 => x"74b00c87",
2297 => x"3d0d04fb",
2298 => x"3d0d800b",
2299 => x"80e0fc0c",
2300 => x"7a537952",
2301 => x"78518299",
2302 => x"3fb00855",
2303 => x"b008ff2e",
2304 => x"883874b0",
2305 => x"0c873d0d",
2306 => x"0480e0fc",
2307 => x"08567580",
2308 => x"2ef03877",
2309 => x"76710c54",
2310 => x"74b00c87",
2311 => x"3d0d04fe",
2312 => x"3d0d80e0",
2313 => x"f0085170",
2314 => x"8a3880e1",
2315 => x"807080e0",
2316 => x"f00c5170",
2317 => x"75125252",
2318 => x"ff537087",
2319 => x"fb808026",
2320 => x"88387080",
2321 => x"e0f00c71",
2322 => x"5372b00c",
2323 => x"843d0d04",
2324 => x"fd3d0d80",
2325 => x"0b80d0f4",
2326 => x"08545472",
2327 => x"812e9c38",
2328 => x"7380e0f4",
2329 => x"0cc0ff3f",
2330 => x"ffbf953f",
2331 => x"80e0c852",
2332 => x"8151c38a",
2333 => x"3fb00851",
2334 => x"85c63f72",
2335 => x"80e0f40c",
2336 => x"c0e43fff",
2337 => x"befa3f80",
2338 => x"e0c85281",
2339 => x"51c2ef3f",
2340 => x"b0085185",
2341 => x"ab3f00ff",
2342 => x"39f53d0d",
2343 => x"7e6080e0",
2344 => x"f408705b",
2345 => x"585b5b75",
2346 => x"80c53877",
2347 => x"7a25a238",
2348 => x"771b7033",
2349 => x"7081ff06",
2350 => x"58585975",
2351 => x"8a2e9938",
2352 => x"7681ff06",
2353 => x"51ffbffd",
2354 => x"3f811858",
2355 => x"797824e0",
2356 => x"3879b00c",
2357 => x"8d3d0d04",
2358 => x"8d51ffbf",
2359 => x"e83f7833",
2360 => x"7081ff06",
2361 => x"5257ffbf",
2362 => x"dc3f8118",
2363 => x"58de3979",
2364 => x"557a547d",
2365 => x"5385528d",
2366 => x"3dfc0551",
2367 => x"ffbec33f",
2368 => x"b0085684",
2369 => x"b43f7bb0",
2370 => x"080c75b0",
2371 => x"0c8d3d0d",
2372 => x"04f63d0d",
2373 => x"7d7f80e0",
2374 => x"f408705b",
2375 => x"585a5a75",
2376 => x"80c43877",
2377 => x"7925b638",
2378 => x"ffbef53f",
2379 => x"b00881ff",
2380 => x"06708d32",
2381 => x"7030709f",
2382 => x"2a515157",
2383 => x"57768a2e",
2384 => x"80c63875",
2385 => x"802e80c0",
2386 => x"38771a56",
2387 => x"76763476",
2388 => x"51ffbef1",
2389 => x"3f811858",
2390 => x"787824cc",
2391 => x"38775675",
2392 => x"b00c8c3d",
2393 => x"0d047855",
2394 => x"79547c53",
2395 => x"84528c3d",
2396 => x"fc0551ff",
2397 => x"bdcc3fb0",
2398 => x"085683bd",
2399 => x"3f7ab008",
2400 => x"0c75b00c",
2401 => x"8c3d0d04",
2402 => x"771a568a",
2403 => x"76348118",
2404 => x"588d51ff",
2405 => x"beaf3f8a",
2406 => x"51ffbea9",
2407 => x"3f7756ff",
2408 => x"be39fb3d",
2409 => x"0d80e0f4",
2410 => x"08705654",
2411 => x"73883874",
2412 => x"b00c873d",
2413 => x"0d047753",
2414 => x"8352873d",
2415 => x"fc0551ff",
2416 => x"bd803fb0",
2417 => x"085482f1",
2418 => x"3f75b008",
2419 => x"0c73b00c",
2420 => x"873d0d04",
2421 => x"fa3d0d80",
2422 => x"e0f40880",
2423 => x"2ea3387a",
2424 => x"55795478",
2425 => x"53865288",
2426 => x"3dfc0551",
2427 => x"ffbcd33f",
2428 => x"b0085682",
2429 => x"c43f76b0",
2430 => x"080c75b0",
2431 => x"0c883d0d",
2432 => x"0482b63f",
2433 => x"9d0bb008",
2434 => x"0cff0bb0",
2435 => x"0c883d0d",
2436 => x"04fb3d0d",
2437 => x"77795656",
2438 => x"80705454",
2439 => x"7375259f",
2440 => x"38741010",
2441 => x"10f80552",
2442 => x"72167033",
2443 => x"70742b76",
2444 => x"078116f8",
2445 => x"16565656",
2446 => x"51517473",
2447 => x"24ea3873",
2448 => x"b00c873d",
2449 => x"0d04fc3d",
2450 => x"0d767855",
2451 => x"55bc5380",
2452 => x"527351f5",
2453 => x"be3f8452",
2454 => x"7451ffb5",
2455 => x"3fb00874",
2456 => x"23845284",
2457 => x"1551ffa9",
2458 => x"3fb00882",
2459 => x"15238452",
2460 => x"881551ff",
2461 => x"9c3fb008",
2462 => x"84150c84",
2463 => x"528c1551",
2464 => x"ff8f3fb0",
2465 => x"08881523",
2466 => x"84529015",
2467 => x"51ff823f",
2468 => x"b0088a15",
2469 => x"23845294",
2470 => x"1551fef5",
2471 => x"3fb0088c",
2472 => x"15238452",
2473 => x"981551fe",
2474 => x"e83fb008",
2475 => x"8e152388",
2476 => x"529c1551",
2477 => x"fedb3fb0",
2478 => x"0890150c",
2479 => x"863d0d04",
2480 => x"e93d0d6a",
2481 => x"80e0f408",
2482 => x"57577593",
2483 => x"3880c080",
2484 => x"0b84180c",
2485 => x"75ac180c",
2486 => x"75b00c99",
2487 => x"3d0d0489",
2488 => x"3d70556a",
2489 => x"54558a52",
2490 => x"993dffbc",
2491 => x"0551ffba",
2492 => x"d13fb008",
2493 => x"77537552",
2494 => x"56fecb3f",
2495 => x"bc3f77b0",
2496 => x"080c75b0",
2497 => x"0c993d0d",
2498 => x"04fc3d0d",
2499 => x"815480e0",
2500 => x"f4088838",
2501 => x"73b00c86",
2502 => x"3d0d0476",
2503 => x"5397b952",
2504 => x"863dfc05",
2505 => x"51ffba9a",
2506 => x"3fb00854",
2507 => x"8c3f74b0",
2508 => x"080c73b0",
2509 => x"0c863d0d",
2510 => x"0480d184",
2511 => x"08b00c04",
2512 => x"f73d0d7b",
2513 => x"80d18408",
2514 => x"82c81108",
2515 => x"5a545a77",
2516 => x"802e80da",
2517 => x"38818818",
2518 => x"841908ff",
2519 => x"0581712b",
2520 => x"59555980",
2521 => x"742480ea",
2522 => x"38807424",
2523 => x"b5387382",
2524 => x"2b781188",
2525 => x"05565681",
2526 => x"80190877",
2527 => x"06537280",
2528 => x"2eb63878",
2529 => x"16700853",
2530 => x"53795174",
2531 => x"0853722d",
2532 => x"ff14fc17",
2533 => x"fc177981",
2534 => x"2c5a5757",
2535 => x"54738025",
2536 => x"d6387708",
2537 => x"5877ffad",
2538 => x"3880d184",
2539 => x"0853bc13",
2540 => x"08a53879",
2541 => x"51f9df3f",
2542 => x"74085372",
2543 => x"2dff14fc",
2544 => x"17fc1779",
2545 => x"812c5a57",
2546 => x"57547380",
2547 => x"25ffa838",
2548 => x"d1398057",
2549 => x"ff933972",
2550 => x"51bc1308",
2551 => x"53722d79",
2552 => x"51f9b33f",
2553 => x"ff3d0d80",
2554 => x"e0d00bfc",
2555 => x"05700852",
2556 => x"5270ff2e",
2557 => x"9138702d",
2558 => x"fc127008",
2559 => x"525270ff",
2560 => x"2e098106",
2561 => x"f138833d",
2562 => x"0d0404ff",
2563 => x"bac33f04",
2564 => x"00ffffff",
2565 => x"ff00ffff",
2566 => x"ffff00ff",
2567 => x"ffffff00",
2568 => x"00000040",
2569 => x"30313233",
2570 => x"34353637",
2571 => x"38396162",
2572 => x"63646566",
2573 => x"00000000",
2574 => x"476f7420",
2575 => x"696e7465",
2576 => x"72727570",
2577 => x"740a0000",
2578 => x"633a0000",
2579 => x"733a0000",
2580 => x"4e6f2069",
2581 => x"6e746572",
2582 => x"72757074",
2583 => x"0a000000",
2584 => x"43000000",
2585 => x"64756d6d",
2586 => x"792e6578",
2587 => x"65000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00003058",
2592 => x"00002824",
2593 => x"00002888",
2594 => x"00000000",
2595 => x"00002af0",
2596 => x"00002b4c",
2597 => x"00002ba8",
2598 => x"00000000",
2599 => x"00000000",
2600 => x"00000000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00002860",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000001",
2637 => x"330eabcd",
2638 => x"1234e66d",
2639 => x"deec0005",
2640 => x"000b0000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000000",
2827 => x"00000000",
2828 => x"00000000",
2829 => x"ffffffff",
2830 => x"00000000",
2831 => x"00020000",
2832 => x"00000000",
2833 => x"00000000",
2834 => x"00002c40",
2835 => x"00002c40",
2836 => x"00002c48",
2837 => x"00002c48",
2838 => x"00002c50",
2839 => x"00002c50",
2840 => x"00002c58",
2841 => x"00002c58",
2842 => x"00002c60",
2843 => x"00002c60",
2844 => x"00002c68",
2845 => x"00002c68",
2846 => x"00002c70",
2847 => x"00002c70",
2848 => x"00002c78",
2849 => x"00002c78",
2850 => x"00002c80",
2851 => x"00002c80",
2852 => x"00002c88",
2853 => x"00002c88",
2854 => x"00002c90",
2855 => x"00002c90",
2856 => x"00002c98",
2857 => x"00002c98",
2858 => x"00002ca0",
2859 => x"00002ca0",
2860 => x"00002ca8",
2861 => x"00002ca8",
2862 => x"00002cb0",
2863 => x"00002cb0",
2864 => x"00002cb8",
2865 => x"00002cb8",
2866 => x"00002cc0",
2867 => x"00002cc0",
2868 => x"00002cc8",
2869 => x"00002cc8",
2870 => x"00002cd0",
2871 => x"00002cd0",
2872 => x"00002cd8",
2873 => x"00002cd8",
2874 => x"00002ce0",
2875 => x"00002ce0",
2876 => x"00002ce8",
2877 => x"00002ce8",
2878 => x"00002cf0",
2879 => x"00002cf0",
2880 => x"00002cf8",
2881 => x"00002cf8",
2882 => x"00002d00",
2883 => x"00002d00",
2884 => x"00002d08",
2885 => x"00002d08",
2886 => x"00002d10",
2887 => x"00002d10",
2888 => x"00002d18",
2889 => x"00002d18",
2890 => x"00002d20",
2891 => x"00002d20",
2892 => x"00002d28",
2893 => x"00002d28",
2894 => x"00002d30",
2895 => x"00002d30",
2896 => x"00002d38",
2897 => x"00002d38",
2898 => x"00002d40",
2899 => x"00002d40",
2900 => x"00002d48",
2901 => x"00002d48",
2902 => x"00002d50",
2903 => x"00002d50",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"00002eb8",
2993 => x"00002eb8",
2994 => x"00002ec0",
2995 => x"00002ec0",
2996 => x"00002ec8",
2997 => x"00002ec8",
2998 => x"00002ed0",
2999 => x"00002ed0",
3000 => x"00002ed8",
3001 => x"00002ed8",
3002 => x"00002ee0",
3003 => x"00002ee0",
3004 => x"00002ee8",
3005 => x"00002ee8",
3006 => x"00002ef0",
3007 => x"00002ef0",
3008 => x"00002ef8",
3009 => x"00002ef8",
3010 => x"00002f00",
3011 => x"00002f00",
3012 => x"00002f08",
3013 => x"00002f08",
3014 => x"00002f10",
3015 => x"00002f10",
3016 => x"00002f18",
3017 => x"00002f18",
3018 => x"00002f20",
3019 => x"00002f20",
3020 => x"00002f28",
3021 => x"00002f28",
3022 => x"00002f30",
3023 => x"00002f30",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"00002fa0",
3051 => x"00002fa0",
3052 => x"00002fa8",
3053 => x"00002fa8",
3054 => x"00002fb0",
3055 => x"00002fb0",
3056 => x"00002fb8",
3057 => x"00002fb8",
3058 => x"00002fc0",
3059 => x"00002fc0",
3060 => x"00002fc8",
3061 => x"00002fc8",
3062 => x"00002fd0",
3063 => x"00002fd0",
3064 => x"00002fd8",
3065 => x"00002fd8",
3066 => x"00002fe0",
3067 => x"00002fe0",
3068 => x"00002fe8",
3069 => x"00002fe8",
3070 => x"00002ff0",
3071 => x"00002ff0",
3072 => x"00002ff8",
3073 => x"00002ff8",
3074 => x"00003000",
3075 => x"00003000",
3076 => x"00003008",
3077 => x"00003008",
3078 => x"00003010",
3079 => x"00003010",
3080 => x"00003018",
3081 => x"00003018",
3082 => x"00003020",
3083 => x"00003020",
3084 => x"00003028",
3085 => x"00003028",
3086 => x"00003030",
3087 => x"00003030",
3088 => x"00003038",
3089 => x"00003038",
3090 => x"00002864",
3091 => x"ffffffff",
3092 => x"00000000",
3093 => x"ffffffff",
3094 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

