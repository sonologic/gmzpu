------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(

0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cfa40c",
3 => x"3a0b0b80",
4 => x"c7970400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"0b0b0b89",
9 => x"90040000",
10 => x"00000000",
11 => x"00000000",
12 => x"00000000",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80ce",
162 => x"d0738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"0b0b0b88",
169 => x"f8040000",
170 => x"00000000",
171 => x"00000000",
172 => x"00000000",
173 => x"00000000",
174 => x"00000000",
175 => x"00000000",
176 => x"0b0b0b88",
177 => x"e0040000",
178 => x"00000000",
179 => x"00000000",
180 => x"00000000",
181 => x"00000000",
182 => x"00000000",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cfa00c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83853f80",
257 => x"c69c3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"b008b408",
281 => x"b8087575",
282 => x"8ec72d50",
283 => x"50b00856",
284 => x"b80cb40c",
285 => x"b00c5104",
286 => x"b008b408",
287 => x"b8087575",
288 => x"8d952d50",
289 => x"50b00856",
290 => x"b80cb40c",
291 => x"b00c5104",
292 => x"b008b408",
293 => x"b8088bb6",
294 => x"2db80cb4",
295 => x"0cb00c04",
296 => x"fe3d0d0b",
297 => x"0b80df94",
298 => x"08538413",
299 => x"0870882a",
300 => x"70810651",
301 => x"52527080",
302 => x"2ef03871",
303 => x"81ff06b0",
304 => x"0c843d0d",
305 => x"04ff3d0d",
306 => x"0b0b80df",
307 => x"94085271",
308 => x"0870882a",
309 => x"81327081",
310 => x"06515151",
311 => x"70f13873",
312 => x"720c833d",
313 => x"0d0480cf",
314 => x"a008802e",
315 => x"a43880cf",
316 => x"a408822e",
317 => x"bd388380",
318 => x"800b0b0b",
319 => x"80df940c",
320 => x"82a0800b",
321 => x"80df980c",
322 => x"8290800b",
323 => x"80df9c0c",
324 => x"04f88080",
325 => x"80a40b0b",
326 => x"0b80df94",
327 => x"0cf88080",
328 => x"82800b80",
329 => x"df980cf8",
330 => x"80808480",
331 => x"0b80df9c",
332 => x"0c0480c0",
333 => x"a8808c0b",
334 => x"0b0b80df",
335 => x"940c80c0",
336 => x"a880940b",
337 => x"80df980c",
338 => x"80cee00b",
339 => x"80df9c0c",
340 => x"04ff3d0d",
341 => x"80dfa033",
342 => x"5170a738",
343 => x"80cfac08",
344 => x"70085252",
345 => x"70802e94",
346 => x"38841280",
347 => x"cfac0c70",
348 => x"2d80cfac",
349 => x"08700852",
350 => x"5270ee38",
351 => x"810b80df",
352 => x"a034833d",
353 => x"0d040480",
354 => x"3d0d0b0b",
355 => x"80df9008",
356 => x"802e8e38",
357 => x"0b0b0b0b",
358 => x"800b802e",
359 => x"09810685",
360 => x"38823d0d",
361 => x"040b0b80",
362 => x"df90510b",
363 => x"0b0bf4d0",
364 => x"3f823d0d",
365 => x"0404ff3d",
366 => x"0d8e8080",
367 => x"0880cfb0",
368 => x"08811180",
369 => x"cfb00c52",
370 => x"52800b8e",
371 => x"80800c71",
372 => x"822a8106",
373 => x"5271802e",
374 => x"8738800b",
375 => x"8e908c0c",
376 => x"833d0d04",
377 => x"f73d0d7b",
378 => x"54870b89",
379 => x"3d80cfb4",
380 => x"08585855",
381 => x"7417748f",
382 => x"06175353",
383 => x"71337334",
384 => x"73842aff",
385 => x"16565474",
386 => x"8025e938",
387 => x"800b8b3d",
388 => x"34765186",
389 => x"d53f8b3d",
390 => x"0d04f73d",
391 => x"0d80cef8",
392 => x"5186c73f",
393 => x"800b8c80",
394 => x"800c868d",
395 => x"a00b8e90",
396 => x"840c9e0b",
397 => x"8e90880c",
398 => x"840b8e80",
399 => x"840c80ce",
400 => x"fc5186a6",
401 => x"3f80cfb0",
402 => x"08893d58",
403 => x"5380cfb0",
404 => x"08527272",
405 => x"2ef73880",
406 => x"cf845186",
407 => x"8d3f80cf",
408 => x"b0085487",
409 => x"0b80cfb4",
410 => x"08575574",
411 => x"17748f06",
412 => x"17535371",
413 => x"33733473",
414 => x"842aff16",
415 => x"56547480",
416 => x"25e93880",
417 => x"0b8b3d34",
418 => x"765185de",
419 => x"3f80cfb0",
420 => x"0853ffb9",
421 => x"39bc0802",
422 => x"bc0cf93d",
423 => x"0d800bbc",
424 => x"08fc050c",
425 => x"bc088805",
426 => x"088025ab",
427 => x"38bc0888",
428 => x"050830bc",
429 => x"0888050c",
430 => x"800bbc08",
431 => x"f4050cbc",
432 => x"08fc0508",
433 => x"8838810b",
434 => x"bc08f405",
435 => x"0cbc08f4",
436 => x"0508bc08",
437 => x"fc050cbc",
438 => x"088c0508",
439 => x"8025ab38",
440 => x"bc088c05",
441 => x"0830bc08",
442 => x"8c050c80",
443 => x"0bbc08f0",
444 => x"050cbc08",
445 => x"fc050888",
446 => x"38810bbc",
447 => x"08f0050c",
448 => x"bc08f005",
449 => x"08bc08fc",
450 => x"050c8053",
451 => x"bc088c05",
452 => x"0852bc08",
453 => x"88050851",
454 => x"81a73fb0",
455 => x"0870bc08",
456 => x"f8050c54",
457 => x"bc08fc05",
458 => x"08802e8c",
459 => x"38bc08f8",
460 => x"050830bc",
461 => x"08f8050c",
462 => x"bc08f805",
463 => x"0870b00c",
464 => x"54893d0d",
465 => x"bc0c04bc",
466 => x"0802bc0c",
467 => x"fb3d0d80",
468 => x"0bbc08fc",
469 => x"050cbc08",
470 => x"88050880",
471 => x"259338bc",
472 => x"08880508",
473 => x"30bc0888",
474 => x"050c810b",
475 => x"bc08fc05",
476 => x"0cbc088c",
477 => x"05088025",
478 => x"8c38bc08",
479 => x"8c050830",
480 => x"bc088c05",
481 => x"0c8153bc",
482 => x"088c0508",
483 => x"52bc0888",
484 => x"050851ad",
485 => x"3fb00870",
486 => x"bc08f805",
487 => x"0c54bc08",
488 => x"fc050880",
489 => x"2e8c38bc",
490 => x"08f80508",
491 => x"30bc08f8",
492 => x"050cbc08",
493 => x"f8050870",
494 => x"b00c5487",
495 => x"3d0dbc0c",
496 => x"04bc0802",
497 => x"bc0cfd3d",
498 => x"0d810bbc",
499 => x"08fc050c",
500 => x"800bbc08",
501 => x"f8050cbc",
502 => x"088c0508",
503 => x"bc088805",
504 => x"0827ac38",
505 => x"bc08fc05",
506 => x"08802ea3",
507 => x"38800bbc",
508 => x"088c0508",
509 => x"249938bc",
510 => x"088c0508",
511 => x"10bc088c",
512 => x"050cbc08",
513 => x"fc050810",
514 => x"bc08fc05",
515 => x"0cc939bc",
516 => x"08fc0508",
517 => x"802e80c9",
518 => x"38bc088c",
519 => x"0508bc08",
520 => x"88050826",
521 => x"a138bc08",
522 => x"880508bc",
523 => x"088c0508",
524 => x"31bc0888",
525 => x"050cbc08",
526 => x"f80508bc",
527 => x"08fc0508",
528 => x"07bc08f8",
529 => x"050cbc08",
530 => x"fc050881",
531 => x"2abc08fc",
532 => x"050cbc08",
533 => x"8c050881",
534 => x"2abc088c",
535 => x"050cffaf",
536 => x"39bc0890",
537 => x"0508802e",
538 => x"8f38bc08",
539 => x"88050870",
540 => x"bc08f405",
541 => x"0c518d39",
542 => x"bc08f805",
543 => x"0870bc08",
544 => x"f4050c51",
545 => x"bc08f405",
546 => x"08b00c85",
547 => x"3d0dbc0c",
548 => x"04fc3d0d",
549 => x"7670797b",
550 => x"55555555",
551 => x"8f72278c",
552 => x"38727507",
553 => x"83065170",
554 => x"802ea738",
555 => x"ff125271",
556 => x"ff2e9838",
557 => x"72708105",
558 => x"54337470",
559 => x"81055634",
560 => x"ff125271",
561 => x"ff2e0981",
562 => x"06ea3874",
563 => x"b00c863d",
564 => x"0d047451",
565 => x"72708405",
566 => x"54087170",
567 => x"8405530c",
568 => x"72708405",
569 => x"54087170",
570 => x"8405530c",
571 => x"72708405",
572 => x"54087170",
573 => x"8405530c",
574 => x"72708405",
575 => x"54087170",
576 => x"8405530c",
577 => x"f0125271",
578 => x"8f26c938",
579 => x"83722795",
580 => x"38727084",
581 => x"05540871",
582 => x"70840553",
583 => x"0cfc1252",
584 => x"718326ed",
585 => x"387054ff",
586 => x"8339f73d",
587 => x"0d7c7052",
588 => x"5380c83f",
589 => x"7254b008",
590 => x"5580cf8c",
591 => x"568157b0",
592 => x"0881055a",
593 => x"8b3de411",
594 => x"59538259",
595 => x"f413527b",
596 => x"88110852",
597 => x"5381833f",
598 => x"b0083070",
599 => x"b008079f",
600 => x"2c8a07b0",
601 => x"0c538b3d",
602 => x"0d04ff3d",
603 => x"0d735280",
604 => x"cfb80851",
605 => x"ffb43f83",
606 => x"3d0d04fd",
607 => x"3d0d7570",
608 => x"71830653",
609 => x"555270b8",
610 => x"38717008",
611 => x"7009f7fb",
612 => x"fdff1206",
613 => x"70f88482",
614 => x"81800651",
615 => x"51525370",
616 => x"9d388413",
617 => x"70087009",
618 => x"f7fbfdff",
619 => x"120670f8",
620 => x"84828180",
621 => x"06515152",
622 => x"5370802e",
623 => x"e5387252",
624 => x"71335170",
625 => x"802e8a38",
626 => x"81127033",
627 => x"525270f8",
628 => x"38717431",
629 => x"b00c853d",
630 => x"0d04f23d",
631 => x"0d606288",
632 => x"11087057",
633 => x"575f5a74",
634 => x"802e818f",
635 => x"388c1a22",
636 => x"70832a81",
637 => x"32708106",
638 => x"51555873",
639 => x"8638901a",
640 => x"08913879",
641 => x"5190a13f",
642 => x"ff54b008",
643 => x"80ed388c",
644 => x"1a22587d",
645 => x"08578078",
646 => x"83ffff06",
647 => x"70812a70",
648 => x"81065156",
649 => x"57557375",
650 => x"2e80d738",
651 => x"74903876",
652 => x"08841808",
653 => x"88195956",
654 => x"5974802e",
655 => x"f2387454",
656 => x"88807527",
657 => x"84388880",
658 => x"54735378",
659 => x"529c1a08",
660 => x"51a41a08",
661 => x"54732d80",
662 => x"0bb00825",
663 => x"82e638b0",
664 => x"081975b0",
665 => x"08317f88",
666 => x"0508b008",
667 => x"31706188",
668 => x"050c5656",
669 => x"5973ffb4",
670 => x"38805473",
671 => x"b00c903d",
672 => x"0d047581",
673 => x"32708106",
674 => x"76415154",
675 => x"73802e81",
676 => x"c1387490",
677 => x"38760884",
678 => x"18088819",
679 => x"59565974",
680 => x"802ef238",
681 => x"881a0878",
682 => x"83ffff06",
683 => x"70892a70",
684 => x"81065156",
685 => x"59567380",
686 => x"2e82fa38",
687 => x"7575278d",
688 => x"3877872a",
689 => x"70810651",
690 => x"547382b5",
691 => x"38747627",
692 => x"83387456",
693 => x"75537852",
694 => x"79085185",
695 => x"823f881a",
696 => x"08763188",
697 => x"1b0c7908",
698 => x"167a0c74",
699 => x"56751975",
700 => x"77317f88",
701 => x"05087831",
702 => x"70618805",
703 => x"0c565659",
704 => x"73802efe",
705 => x"f4388c1a",
706 => x"2258ff86",
707 => x"39777854",
708 => x"79537b52",
709 => x"5684c83f",
710 => x"881a0878",
711 => x"31881b0c",
712 => x"7908187a",
713 => x"0c7c7631",
714 => x"5d7c8e38",
715 => x"79518fdb",
716 => x"3fb00881",
717 => x"8f38b008",
718 => x"5f751975",
719 => x"77317f88",
720 => x"05087831",
721 => x"70618805",
722 => x"0c565659",
723 => x"73802efe",
724 => x"a8387481",
725 => x"83387608",
726 => x"84180888",
727 => x"19595659",
728 => x"74802ef2",
729 => x"3874538a",
730 => x"52785182",
731 => x"d33fb008",
732 => x"79318105",
733 => x"5db00884",
734 => x"3881155d",
735 => x"815f7c58",
736 => x"747d2783",
737 => x"38745894",
738 => x"1a08881b",
739 => x"0811575c",
740 => x"807a085c",
741 => x"54901a08",
742 => x"7b278338",
743 => x"81547578",
744 => x"25843873",
745 => x"ba387b78",
746 => x"24fee238",
747 => x"7b537852",
748 => x"9c1a0851",
749 => x"a41a0854",
750 => x"732db008",
751 => x"56b00880",
752 => x"24fee238",
753 => x"8c1a2280",
754 => x"c0075473",
755 => x"8c1b23ff",
756 => x"5473b00c",
757 => x"903d0d04",
758 => x"7effa338",
759 => x"ff873975",
760 => x"5378527a",
761 => x"5182f83f",
762 => x"7908167a",
763 => x"0c79518e",
764 => x"9a3fb008",
765 => x"cf387c76",
766 => x"315d7cfe",
767 => x"bc38feac",
768 => x"39901a08",
769 => x"7a087131",
770 => x"76117056",
771 => x"5a575280",
772 => x"cfb80851",
773 => x"848c3fb0",
774 => x"08802eff",
775 => x"a738b008",
776 => x"901b0cb0",
777 => x"08167a0c",
778 => x"77941b0c",
779 => x"74881b0c",
780 => x"7456fd99",
781 => x"39790858",
782 => x"901a0878",
783 => x"27833881",
784 => x"54757527",
785 => x"843873b3",
786 => x"38941a08",
787 => x"56757526",
788 => x"80d33875",
789 => x"5378529c",
790 => x"1a0851a4",
791 => x"1a085473",
792 => x"2db00856",
793 => x"b0088024",
794 => x"fd83388c",
795 => x"1a2280c0",
796 => x"0754738c",
797 => x"1b23ff54",
798 => x"fed73975",
799 => x"53785277",
800 => x"5181dc3f",
801 => x"7908167a",
802 => x"0c79518c",
803 => x"fe3fb008",
804 => x"802efcd9",
805 => x"388c1a22",
806 => x"80c00754",
807 => x"738c1b23",
808 => x"ff54fead",
809 => x"39747554",
810 => x"79537852",
811 => x"5681b03f",
812 => x"881a0875",
813 => x"31881b0c",
814 => x"7908157a",
815 => x"0cfcae39",
816 => x"fa3d0d7a",
817 => x"79028805",
818 => x"a7053356",
819 => x"52538373",
820 => x"278a3870",
821 => x"83065271",
822 => x"802ea838",
823 => x"ff135372",
824 => x"ff2e9738",
825 => x"70335273",
826 => x"722e9138",
827 => x"8111ff14",
828 => x"545172ff",
829 => x"2e098106",
830 => x"eb388051",
831 => x"70b00c88",
832 => x"3d0d0470",
833 => x"72575583",
834 => x"51758280",
835 => x"2914ff12",
836 => x"52567080",
837 => x"25f33883",
838 => x"7327bf38",
839 => x"74087632",
840 => x"7009f7fb",
841 => x"fdff1206",
842 => x"70f88482",
843 => x"81800651",
844 => x"51517080",
845 => x"2e993874",
846 => x"51805270",
847 => x"33577377",
848 => x"2effb938",
849 => x"81118113",
850 => x"53518372",
851 => x"27ed38fc",
852 => x"13841656",
853 => x"53728326",
854 => x"c3387451",
855 => x"fefe39fa",
856 => x"3d0d787a",
857 => x"7c727272",
858 => x"57575759",
859 => x"56567476",
860 => x"27b23876",
861 => x"15517571",
862 => x"27aa3870",
863 => x"7717ff14",
864 => x"54555371",
865 => x"ff2e9638",
866 => x"ff14ff14",
867 => x"54547233",
868 => x"7434ff12",
869 => x"5271ff2e",
870 => x"098106ec",
871 => x"3875b00c",
872 => x"883d0d04",
873 => x"768f2697",
874 => x"38ff1252",
875 => x"71ff2eed",
876 => x"38727081",
877 => x"05543374",
878 => x"70810556",
879 => x"34eb3974",
880 => x"76078306",
881 => x"5170e238",
882 => x"75755451",
883 => x"72708405",
884 => x"54087170",
885 => x"8405530c",
886 => x"72708405",
887 => x"54087170",
888 => x"8405530c",
889 => x"72708405",
890 => x"54087170",
891 => x"8405530c",
892 => x"72708405",
893 => x"54087170",
894 => x"8405530c",
895 => x"f0125271",
896 => x"8f26c938",
897 => x"83722795",
898 => x"38727084",
899 => x"05540871",
900 => x"70840553",
901 => x"0cfc1252",
902 => x"718326ed",
903 => x"387054ff",
904 => x"8839ef3d",
905 => x"0d636567",
906 => x"405d427b",
907 => x"802e84fa",
908 => x"386151a5",
909 => x"b43ff81c",
910 => x"70841208",
911 => x"70fc0670",
912 => x"628b0570",
913 => x"f8064159",
914 => x"455b5c41",
915 => x"57967427",
916 => x"82c33880",
917 => x"7b247e7c",
918 => x"26075980",
919 => x"5478742e",
920 => x"09810682",
921 => x"a938777b",
922 => x"2581fc38",
923 => x"771780d6",
924 => x"f40b8805",
925 => x"085e567c",
926 => x"762e84bd",
927 => x"38841608",
928 => x"70fe0617",
929 => x"84110881",
930 => x"06515555",
931 => x"73828b38",
932 => x"74fc0659",
933 => x"7c762e84",
934 => x"dd387719",
935 => x"5f7e7b25",
936 => x"81fd3879",
937 => x"81065473",
938 => x"82bf3876",
939 => x"77083184",
940 => x"1108fc06",
941 => x"565a7580",
942 => x"2e91387c",
943 => x"762e84ea",
944 => x"38741918",
945 => x"59787b25",
946 => x"84893879",
947 => x"802e8299",
948 => x"38771556",
949 => x"7a762482",
950 => x"90388c1a",
951 => x"08881b08",
952 => x"718c120c",
953 => x"88120c55",
954 => x"79765957",
955 => x"881761fc",
956 => x"05575975",
957 => x"a42685ef",
958 => x"387b7955",
959 => x"55937627",
960 => x"80c9387b",
961 => x"7084055d",
962 => x"087c5679",
963 => x"0c747084",
964 => x"0556088c",
965 => x"180c9017",
966 => x"549b7627",
967 => x"ae387470",
968 => x"84055608",
969 => x"740c7470",
970 => x"84055608",
971 => x"94180c98",
972 => x"1754a376",
973 => x"27953874",
974 => x"70840556",
975 => x"08740c74",
976 => x"70840556",
977 => x"089c180c",
978 => x"a0175474",
979 => x"70840556",
980 => x"08747084",
981 => x"05560c74",
982 => x"70840556",
983 => x"08747084",
984 => x"05560c74",
985 => x"08740c77",
986 => x"7b315675",
987 => x"8f2680c9",
988 => x"38841708",
989 => x"81067807",
990 => x"84180c77",
991 => x"17841108",
992 => x"81078412",
993 => x"0c546151",
994 => x"a2e03f88",
995 => x"175473b0",
996 => x"0c933d0d",
997 => x"04905bfd",
998 => x"ba397856",
999 => x"fe85398c",
1000 => x"16088817",
1001 => x"08718c12",
1002 => x"0c88120c",
1003 => x"557e707c",
1004 => x"3157588f",
1005 => x"7627ffb9",
1006 => x"387a1784",
1007 => x"18088106",
1008 => x"7c078419",
1009 => x"0c768107",
1010 => x"84120c76",
1011 => x"11841108",
1012 => x"81078412",
1013 => x"0c558805",
1014 => x"5261518c",
1015 => x"f63f6151",
1016 => x"a2883f88",
1017 => x"1754ffa6",
1018 => x"397d5261",
1019 => x"5194f53f",
1020 => x"b00859b0",
1021 => x"08802e81",
1022 => x"a338b008",
1023 => x"f8056084",
1024 => x"0508fe06",
1025 => x"61055557",
1026 => x"76742e83",
1027 => x"e638fc18",
1028 => x"5675a426",
1029 => x"81aa387b",
1030 => x"b0085555",
1031 => x"93762780",
1032 => x"d8387470",
1033 => x"84055608",
1034 => x"b0087084",
1035 => x"05b00c0c",
1036 => x"b0087570",
1037 => x"84055708",
1038 => x"71708405",
1039 => x"530c549b",
1040 => x"7627b638",
1041 => x"74708405",
1042 => x"56087470",
1043 => x"8405560c",
1044 => x"74708405",
1045 => x"56087470",
1046 => x"8405560c",
1047 => x"a3762799",
1048 => x"38747084",
1049 => x"05560874",
1050 => x"70840556",
1051 => x"0c747084",
1052 => x"05560874",
1053 => x"70840556",
1054 => x"0c747084",
1055 => x"05560874",
1056 => x"70840556",
1057 => x"0c747084",
1058 => x"05560874",
1059 => x"70840556",
1060 => x"0c740874",
1061 => x"0c7b5261",
1062 => x"518bb83f",
1063 => x"6151a0ca",
1064 => x"3f785473",
1065 => x"b00c933d",
1066 => x"0d047d52",
1067 => x"615193b4",
1068 => x"3fb008b0",
1069 => x"0c933d0d",
1070 => x"04841608",
1071 => x"55fbd139",
1072 => x"75537b52",
1073 => x"b00851ef",
1074 => x"c83f7b52",
1075 => x"61518b83",
1076 => x"3fca398c",
1077 => x"16088817",
1078 => x"08718c12",
1079 => x"0c88120c",
1080 => x"558c1a08",
1081 => x"881b0871",
1082 => x"8c120c88",
1083 => x"120c5579",
1084 => x"795957fb",
1085 => x"f7397719",
1086 => x"901c5555",
1087 => x"737524fb",
1088 => x"a2387a17",
1089 => x"7080d6f4",
1090 => x"0b88050c",
1091 => x"757c3181",
1092 => x"0784120c",
1093 => x"5d841708",
1094 => x"81067b07",
1095 => x"84180c61",
1096 => x"519fc73f",
1097 => x"881754fc",
1098 => x"e5397419",
1099 => x"18901c55",
1100 => x"5d737d24",
1101 => x"fb95388c",
1102 => x"1a08881b",
1103 => x"08718c12",
1104 => x"0c88120c",
1105 => x"55881a61",
1106 => x"fc055759",
1107 => x"75a42681",
1108 => x"ae387b79",
1109 => x"55559376",
1110 => x"2780c938",
1111 => x"7b708405",
1112 => x"5d087c56",
1113 => x"790c7470",
1114 => x"84055608",
1115 => x"8c1b0c90",
1116 => x"1a549b76",
1117 => x"27ae3874",
1118 => x"70840556",
1119 => x"08740c74",
1120 => x"70840556",
1121 => x"08941b0c",
1122 => x"981a54a3",
1123 => x"76279538",
1124 => x"74708405",
1125 => x"5608740c",
1126 => x"74708405",
1127 => x"56089c1b",
1128 => x"0ca01a54",
1129 => x"74708405",
1130 => x"56087470",
1131 => x"8405560c",
1132 => x"74708405",
1133 => x"56087470",
1134 => x"8405560c",
1135 => x"7408740c",
1136 => x"7a1a7080",
1137 => x"d6f40b88",
1138 => x"050c7d7c",
1139 => x"31810784",
1140 => x"120c5484",
1141 => x"1a088106",
1142 => x"7b07841b",
1143 => x"0c61519e",
1144 => x"893f7854",
1145 => x"fdbd3975",
1146 => x"537b5278",
1147 => x"51eda23f",
1148 => x"faf53984",
1149 => x"1708fc06",
1150 => x"18605858",
1151 => x"fae93975",
1152 => x"537b5278",
1153 => x"51ed8a3f",
1154 => x"7a1a7080",
1155 => x"d6f40b88",
1156 => x"050c7d7c",
1157 => x"31810784",
1158 => x"120c5484",
1159 => x"1a088106",
1160 => x"7b07841b",
1161 => x"0cffb639",
1162 => x"fa3d0d78",
1163 => x"80cfb808",
1164 => x"5455b813",
1165 => x"08802e81",
1166 => x"b5388c15",
1167 => x"227083ff",
1168 => x"ff067083",
1169 => x"2a813270",
1170 => x"81065155",
1171 => x"55567280",
1172 => x"2e80dc38",
1173 => x"73842a81",
1174 => x"32810657",
1175 => x"ff537680",
1176 => x"f6387382",
1177 => x"2a708106",
1178 => x"51537280",
1179 => x"2eb938b0",
1180 => x"15085473",
1181 => x"802e9c38",
1182 => x"80c01553",
1183 => x"73732e8f",
1184 => x"38735280",
1185 => x"cfb80851",
1186 => x"87c93f8c",
1187 => x"15225676",
1188 => x"b0160c75",
1189 => x"db065372",
1190 => x"8c162380",
1191 => x"0b84160c",
1192 => x"90150875",
1193 => x"0c725675",
1194 => x"88075372",
1195 => x"8c162390",
1196 => x"1508802e",
1197 => x"80c0388c",
1198 => x"15227081",
1199 => x"06555373",
1200 => x"9d387281",
1201 => x"2a708106",
1202 => x"51537285",
1203 => x"38941508",
1204 => x"54738816",
1205 => x"0c805372",
1206 => x"b00c883d",
1207 => x"0d04800b",
1208 => x"88160c94",
1209 => x"15083098",
1210 => x"160c8053",
1211 => x"ea397251",
1212 => x"82fb3ffe",
1213 => x"c5397451",
1214 => x"8ce83f8c",
1215 => x"15227081",
1216 => x"06555373",
1217 => x"802effba",
1218 => x"38d439f8",
1219 => x"3d0d7a58",
1220 => x"77802e81",
1221 => x"993880cf",
1222 => x"b80854b8",
1223 => x"1408802e",
1224 => x"80ed388c",
1225 => x"18227090",
1226 => x"2b70902c",
1227 => x"70832a81",
1228 => x"3281065c",
1229 => x"51575478",
1230 => x"80cd3890",
1231 => x"18085776",
1232 => x"802e80c3",
1233 => x"38770877",
1234 => x"3177790c",
1235 => x"7683067a",
1236 => x"58555573",
1237 => x"85389418",
1238 => x"08567588",
1239 => x"190c8075",
1240 => x"25a53874",
1241 => x"5376529c",
1242 => x"180851a4",
1243 => x"18085473",
1244 => x"2d800bb0",
1245 => x"082580c9",
1246 => x"38b00817",
1247 => x"75b00831",
1248 => x"56577480",
1249 => x"24dd3880",
1250 => x"0bb00c8a",
1251 => x"3d0d0473",
1252 => x"5181da3f",
1253 => x"8c182270",
1254 => x"902b7090",
1255 => x"2c70832a",
1256 => x"81328106",
1257 => x"5c515754",
1258 => x"78dd38ff",
1259 => x"8e39a68b",
1260 => x"5280cfb8",
1261 => x"085189f1",
1262 => x"3fb008b0",
1263 => x"0c8a3d0d",
1264 => x"048c1822",
1265 => x"80c00754",
1266 => x"738c1923",
1267 => x"ff0bb00c",
1268 => x"8a3d0d04",
1269 => x"803d0d72",
1270 => x"5180710c",
1271 => x"800b8412",
1272 => x"0c800b88",
1273 => x"120c028e",
1274 => x"05228c12",
1275 => x"23029205",
1276 => x"228e1223",
1277 => x"800b9012",
1278 => x"0c800b94",
1279 => x"120c800b",
1280 => x"98120c70",
1281 => x"9c120c80",
1282 => x"c29f0ba0",
1283 => x"120c80c2",
1284 => x"eb0ba412",
1285 => x"0c80c3e7",
1286 => x"0ba8120c",
1287 => x"80c4b80b",
1288 => x"ac120c82",
1289 => x"3d0d04fa",
1290 => x"3d0d7970",
1291 => x"80dc298c",
1292 => x"11547a53",
1293 => x"56578cac",
1294 => x"3fb008b0",
1295 => x"085556b0",
1296 => x"08802ea2",
1297 => x"38b0088c",
1298 => x"0554800b",
1299 => x"b0080c76",
1300 => x"b0088405",
1301 => x"0c73b008",
1302 => x"88050c74",
1303 => x"53805273",
1304 => x"5197f73f",
1305 => x"755473b0",
1306 => x"0c883d0d",
1307 => x"04fc3d0d",
1308 => x"76ab800b",
1309 => x"bc120c55",
1310 => x"810bb816",
1311 => x"0c800b84",
1312 => x"dc160c83",
1313 => x"0b84e016",
1314 => x"0c84e815",
1315 => x"84e4160c",
1316 => x"74548053",
1317 => x"84528415",
1318 => x"0851feb8",
1319 => x"3f745481",
1320 => x"53895288",
1321 => x"150851fe",
1322 => x"ab3f7454",
1323 => x"82538a52",
1324 => x"8c150851",
1325 => x"fe9e3f86",
1326 => x"3d0d04f9",
1327 => x"3d0d7980",
1328 => x"cfb80854",
1329 => x"57b81308",
1330 => x"802e80c8",
1331 => x"3884dc13",
1332 => x"56881608",
1333 => x"841708ff",
1334 => x"05555580",
1335 => x"74249f38",
1336 => x"8c152270",
1337 => x"902b7090",
1338 => x"2c515458",
1339 => x"72802e80",
1340 => x"ca3880dc",
1341 => x"15ff1555",
1342 => x"55738025",
1343 => x"e3387508",
1344 => x"5372802e",
1345 => x"9f387256",
1346 => x"88160884",
1347 => x"1708ff05",
1348 => x"5555c839",
1349 => x"7251fed5",
1350 => x"3f80cfb8",
1351 => x"0884dc05",
1352 => x"56ffae39",
1353 => x"84527651",
1354 => x"fdfd3fb0",
1355 => x"08760cb0",
1356 => x"08802e80",
1357 => x"c038b008",
1358 => x"56ce3981",
1359 => x"0b8c1623",
1360 => x"72750c72",
1361 => x"88160c72",
1362 => x"84160c72",
1363 => x"90160c72",
1364 => x"94160c72",
1365 => x"98160cff",
1366 => x"0b8e1623",
1367 => x"72b0160c",
1368 => x"72b4160c",
1369 => x"7280c416",
1370 => x"0c7280c8",
1371 => x"160c74b0",
1372 => x"0c893d0d",
1373 => x"048c770c",
1374 => x"800bb00c",
1375 => x"893d0d04",
1376 => x"ff3d0da6",
1377 => x"8b527351",
1378 => x"869f3f83",
1379 => x"3d0d0480",
1380 => x"3d0d80cf",
1381 => x"b80851e8",
1382 => x"3f823d0d",
1383 => x"04fb3d0d",
1384 => x"77705256",
1385 => x"96c33f80",
1386 => x"d6f40b88",
1387 => x"05088411",
1388 => x"08fc0670",
1389 => x"7b319fef",
1390 => x"05e08006",
1391 => x"e0800556",
1392 => x"5653a080",
1393 => x"74249438",
1394 => x"80527551",
1395 => x"969d3f80",
1396 => x"d6fc0815",
1397 => x"5372b008",
1398 => x"2e8f3875",
1399 => x"51968b3f",
1400 => x"805372b0",
1401 => x"0c873d0d",
1402 => x"04733052",
1403 => x"755195fb",
1404 => x"3fb008ff",
1405 => x"2ea83880",
1406 => x"d6f40b88",
1407 => x"05087575",
1408 => x"31810784",
1409 => x"120c5380",
1410 => x"d6b80874",
1411 => x"3180d6b8",
1412 => x"0c755195",
1413 => x"d53f810b",
1414 => x"b00c873d",
1415 => x"0d048052",
1416 => x"755195c7",
1417 => x"3f80d6f4",
1418 => x"0b880508",
1419 => x"b0087131",
1420 => x"56538f75",
1421 => x"25ffa438",
1422 => x"b00880d6",
1423 => x"e8083180",
1424 => x"d6b80c74",
1425 => x"81078414",
1426 => x"0c755195",
1427 => x"9d3f8053",
1428 => x"ff9039f6",
1429 => x"3d0d7c7e",
1430 => x"545b7280",
1431 => x"2e828338",
1432 => x"7a519585",
1433 => x"3ff81384",
1434 => x"110870fe",
1435 => x"06701384",
1436 => x"1108fc06",
1437 => x"5d585954",
1438 => x"5880d6fc",
1439 => x"08752e82",
1440 => x"de387884",
1441 => x"160c8073",
1442 => x"8106545a",
1443 => x"727a2e81",
1444 => x"d5387815",
1445 => x"84110881",
1446 => x"06515372",
1447 => x"a0387817",
1448 => x"577981e6",
1449 => x"38881508",
1450 => x"537280d6",
1451 => x"fc2e82f9",
1452 => x"388c1508",
1453 => x"708c150c",
1454 => x"7388120c",
1455 => x"56768107",
1456 => x"84190c76",
1457 => x"1877710c",
1458 => x"53798191",
1459 => x"3883ff77",
1460 => x"2781c838",
1461 => x"76892a77",
1462 => x"832a5653",
1463 => x"72802ebf",
1464 => x"3876862a",
1465 => x"b8055584",
1466 => x"7327b438",
1467 => x"80db1355",
1468 => x"947327ab",
1469 => x"38768c2a",
1470 => x"80ee0555",
1471 => x"80d47327",
1472 => x"9e38768f",
1473 => x"2a80f705",
1474 => x"5582d473",
1475 => x"27913876",
1476 => x"922a80fc",
1477 => x"05558ad4",
1478 => x"73278438",
1479 => x"80fe5574",
1480 => x"10101080",
1481 => x"d6f40588",
1482 => x"11085556",
1483 => x"73762e82",
1484 => x"b3388414",
1485 => x"08fc0653",
1486 => x"7673278d",
1487 => x"38881408",
1488 => x"5473762e",
1489 => x"098106ea",
1490 => x"388c1408",
1491 => x"708c1a0c",
1492 => x"74881a0c",
1493 => x"7888120c",
1494 => x"56778c15",
1495 => x"0c7a5193",
1496 => x"893f8c3d",
1497 => x"0d047708",
1498 => x"78713159",
1499 => x"77058819",
1500 => x"08545772",
1501 => x"80d6fc2e",
1502 => x"80e0388c",
1503 => x"1808708c",
1504 => x"150c7388",
1505 => x"120c56fe",
1506 => x"89398815",
1507 => x"088c1608",
1508 => x"708c130c",
1509 => x"5788170c",
1510 => x"fea33976",
1511 => x"832a7054",
1512 => x"55807524",
1513 => x"81983872",
1514 => x"822c8171",
1515 => x"2b80d6f8",
1516 => x"080780d6",
1517 => x"f40b8405",
1518 => x"0c537410",
1519 => x"101080d6",
1520 => x"f4058811",
1521 => x"08555675",
1522 => x"8c190c73",
1523 => x"88190c77",
1524 => x"88170c77",
1525 => x"8c150cff",
1526 => x"8439815a",
1527 => x"fdb43978",
1528 => x"17738106",
1529 => x"54577298",
1530 => x"38770878",
1531 => x"71315977",
1532 => x"058c1908",
1533 => x"881a0871",
1534 => x"8c120c88",
1535 => x"120c5757",
1536 => x"76810784",
1537 => x"190c7780",
1538 => x"d6f40b88",
1539 => x"050c80d6",
1540 => x"f0087726",
1541 => x"fec73880",
1542 => x"d6ec0852",
1543 => x"7a51fafd",
1544 => x"3f7a5191",
1545 => x"c53ffeba",
1546 => x"3981788c",
1547 => x"150c7888",
1548 => x"150c738c",
1549 => x"1a0c7388",
1550 => x"1a0c5afd",
1551 => x"80398315",
1552 => x"70822c81",
1553 => x"712b80d6",
1554 => x"f8080780",
1555 => x"d6f40b84",
1556 => x"050c5153",
1557 => x"74101010",
1558 => x"80d6f405",
1559 => x"88110855",
1560 => x"56fee439",
1561 => x"74538075",
1562 => x"24a73872",
1563 => x"822c8171",
1564 => x"2b80d6f8",
1565 => x"080780d6",
1566 => x"f40b8405",
1567 => x"0c53758c",
1568 => x"190c7388",
1569 => x"190c7788",
1570 => x"170c778c",
1571 => x"150cfdcd",
1572 => x"39831570",
1573 => x"822c8171",
1574 => x"2b80d6f8",
1575 => x"080780d6",
1576 => x"f40b8405",
1577 => x"0c5153d6",
1578 => x"39f93d0d",
1579 => x"797b5853",
1580 => x"800b80cf",
1581 => x"b8085356",
1582 => x"72722e80",
1583 => x"c03884dc",
1584 => x"13557476",
1585 => x"2eb73888",
1586 => x"15088416",
1587 => x"08ff0554",
1588 => x"54807324",
1589 => x"9d388c14",
1590 => x"2270902b",
1591 => x"70902c51",
1592 => x"53587180",
1593 => x"d83880dc",
1594 => x"14ff1454",
1595 => x"54728025",
1596 => x"e5387408",
1597 => x"5574d038",
1598 => x"80cfb808",
1599 => x"5284dc12",
1600 => x"5574802e",
1601 => x"b1388815",
1602 => x"08841608",
1603 => x"ff055454",
1604 => x"8073249c",
1605 => x"388c1422",
1606 => x"70902b70",
1607 => x"902c5153",
1608 => x"5871ad38",
1609 => x"80dc14ff",
1610 => x"14545472",
1611 => x"8025e638",
1612 => x"74085574",
1613 => x"d13875b0",
1614 => x"0c893d0d",
1615 => x"04735176",
1616 => x"2d75b008",
1617 => x"0780dc15",
1618 => x"ff155555",
1619 => x"56ff9e39",
1620 => x"7351762d",
1621 => x"75b00807",
1622 => x"80dc15ff",
1623 => x"15555556",
1624 => x"ca39ea3d",
1625 => x"0d688c11",
1626 => x"2270812a",
1627 => x"81065758",
1628 => x"567480e4",
1629 => x"388e1622",
1630 => x"70902b70",
1631 => x"902c5155",
1632 => x"58807424",
1633 => x"b138983d",
1634 => x"c4055373",
1635 => x"5280cfb8",
1636 => x"085192ac",
1637 => x"3f800bb0",
1638 => x"08249738",
1639 => x"7983e080",
1640 => x"06547380",
1641 => x"c0802e81",
1642 => x"8f387382",
1643 => x"80802e81",
1644 => x"91388c16",
1645 => x"22577690",
1646 => x"80075473",
1647 => x"8c172388",
1648 => x"805280cf",
1649 => x"b8085181",
1650 => x"9b3fb008",
1651 => x"9d388c16",
1652 => x"22820754",
1653 => x"738c1723",
1654 => x"80c31670",
1655 => x"770c9017",
1656 => x"0c810b94",
1657 => x"170c983d",
1658 => x"0d0480cf",
1659 => x"b808ab80",
1660 => x"0bbc120c",
1661 => x"548c1622",
1662 => x"81800754",
1663 => x"738c1723",
1664 => x"b008760c",
1665 => x"b0089017",
1666 => x"0c88800b",
1667 => x"94170c74",
1668 => x"802ed338",
1669 => x"8e162270",
1670 => x"902b7090",
1671 => x"2c535558",
1672 => x"98a53fb0",
1673 => x"08802eff",
1674 => x"bd388c16",
1675 => x"22810754",
1676 => x"738c1723",
1677 => x"983d0d04",
1678 => x"810b8c17",
1679 => x"225855fe",
1680 => x"f539a816",
1681 => x"0880c3e7",
1682 => x"2e098106",
1683 => x"fee4388c",
1684 => x"16228880",
1685 => x"0754738c",
1686 => x"17238880",
1687 => x"0b80cc17",
1688 => x"0cfedc39",
1689 => x"f33d0d7f",
1690 => x"618b1170",
1691 => x"f8065c55",
1692 => x"555e7296",
1693 => x"26833890",
1694 => x"59807924",
1695 => x"747a2607",
1696 => x"53805472",
1697 => x"742e0981",
1698 => x"0680cb38",
1699 => x"7d518cd9",
1700 => x"3f7883f7",
1701 => x"2680c638",
1702 => x"78832a70",
1703 => x"10101080",
1704 => x"d6f4058c",
1705 => x"11085959",
1706 => x"5a76782e",
1707 => x"83b03884",
1708 => x"1708fc06",
1709 => x"568c1708",
1710 => x"88180871",
1711 => x"8c120c88",
1712 => x"120c5875",
1713 => x"17841108",
1714 => x"81078412",
1715 => x"0c537d51",
1716 => x"8c983f88",
1717 => x"175473b0",
1718 => x"0c8f3d0d",
1719 => x"0478892a",
1720 => x"79832a5b",
1721 => x"5372802e",
1722 => x"bf387886",
1723 => x"2ab8055a",
1724 => x"847327b4",
1725 => x"3880db13",
1726 => x"5a947327",
1727 => x"ab38788c",
1728 => x"2a80ee05",
1729 => x"5a80d473",
1730 => x"279e3878",
1731 => x"8f2a80f7",
1732 => x"055a82d4",
1733 => x"73279138",
1734 => x"78922a80",
1735 => x"fc055a8a",
1736 => x"d4732784",
1737 => x"3880fe5a",
1738 => x"79101010",
1739 => x"80d6f405",
1740 => x"8c110858",
1741 => x"5576752e",
1742 => x"a3388417",
1743 => x"08fc0670",
1744 => x"7a315556",
1745 => x"738f2488",
1746 => x"d5387380",
1747 => x"25fee638",
1748 => x"8c170857",
1749 => x"76752e09",
1750 => x"8106df38",
1751 => x"811a5a80",
1752 => x"d7840857",
1753 => x"7680d6fc",
1754 => x"2e82c038",
1755 => x"841708fc",
1756 => x"06707a31",
1757 => x"5556738f",
1758 => x"2481f938",
1759 => x"80d6fc0b",
1760 => x"80d7880c",
1761 => x"80d6fc0b",
1762 => x"80d7840c",
1763 => x"738025fe",
1764 => x"b23883ff",
1765 => x"762783df",
1766 => x"3875892a",
1767 => x"76832a55",
1768 => x"5372802e",
1769 => x"bf387586",
1770 => x"2ab80554",
1771 => x"847327b4",
1772 => x"3880db13",
1773 => x"54947327",
1774 => x"ab38758c",
1775 => x"2a80ee05",
1776 => x"5480d473",
1777 => x"279e3875",
1778 => x"8f2a80f7",
1779 => x"055482d4",
1780 => x"73279138",
1781 => x"75922a80",
1782 => x"fc05548a",
1783 => x"d4732784",
1784 => x"3880fe54",
1785 => x"73101010",
1786 => x"80d6f405",
1787 => x"88110856",
1788 => x"5874782e",
1789 => x"86cf3884",
1790 => x"1508fc06",
1791 => x"53757327",
1792 => x"8d388815",
1793 => x"08557478",
1794 => x"2e098106",
1795 => x"ea388c15",
1796 => x"0880d6f4",
1797 => x"0b840508",
1798 => x"718c1a0c",
1799 => x"76881a0c",
1800 => x"7888130c",
1801 => x"788c180c",
1802 => x"5d587953",
1803 => x"807a2483",
1804 => x"e6387282",
1805 => x"2c81712b",
1806 => x"5c537a7c",
1807 => x"26819838",
1808 => x"7b7b0653",
1809 => x"7282f138",
1810 => x"79fc0684",
1811 => x"055a7a10",
1812 => x"707d0654",
1813 => x"5b7282e0",
1814 => x"38841a5a",
1815 => x"f1398817",
1816 => x"8c110858",
1817 => x"5876782e",
1818 => x"098106fc",
1819 => x"c238821a",
1820 => x"5afdec39",
1821 => x"78177981",
1822 => x"0784190c",
1823 => x"7080d788",
1824 => x"0c7080d7",
1825 => x"840c80d6",
1826 => x"fc0b8c12",
1827 => x"0c8c1108",
1828 => x"88120c74",
1829 => x"81078412",
1830 => x"0c741175",
1831 => x"710c5153",
1832 => x"7d5188c6",
1833 => x"3f881754",
1834 => x"fcac3980",
1835 => x"d6f40b84",
1836 => x"05087a54",
1837 => x"5c798025",
1838 => x"fef83882",
1839 => x"da397a09",
1840 => x"7c067080",
1841 => x"d6f40b84",
1842 => x"050c5c7a",
1843 => x"105b7a7c",
1844 => x"2685387a",
1845 => x"85b83880",
1846 => x"d6f40b88",
1847 => x"05087084",
1848 => x"1208fc06",
1849 => x"707c317c",
1850 => x"72268f72",
1851 => x"25075757",
1852 => x"5c5d5572",
1853 => x"802e80db",
1854 => x"38797a16",
1855 => x"80d6ec08",
1856 => x"1b90115a",
1857 => x"55575b80",
1858 => x"d6e808ff",
1859 => x"2e8838a0",
1860 => x"8f13e080",
1861 => x"06577652",
1862 => x"7d5187cf",
1863 => x"3fb00854",
1864 => x"b008ff2e",
1865 => x"9038b008",
1866 => x"76278299",
1867 => x"387480d6",
1868 => x"f42e8291",
1869 => x"3880d6f4",
1870 => x"0b880508",
1871 => x"55841508",
1872 => x"fc06707a",
1873 => x"317a7226",
1874 => x"8f722507",
1875 => x"52555372",
1876 => x"83e63874",
1877 => x"79810784",
1878 => x"170c7916",
1879 => x"7080d6f4",
1880 => x"0b88050c",
1881 => x"75810784",
1882 => x"120c547e",
1883 => x"525786fa",
1884 => x"3f881754",
1885 => x"fae03975",
1886 => x"832a7054",
1887 => x"54807424",
1888 => x"819b3872",
1889 => x"822c8171",
1890 => x"2b80d6f8",
1891 => x"08077080",
1892 => x"d6f40b84",
1893 => x"050c7510",
1894 => x"101080d6",
1895 => x"f4058811",
1896 => x"08585a5d",
1897 => x"53778c18",
1898 => x"0c748818",
1899 => x"0c768819",
1900 => x"0c768c16",
1901 => x"0cfcf339",
1902 => x"797a1010",
1903 => x"1080d6f4",
1904 => x"05705759",
1905 => x"5d8c1508",
1906 => x"5776752e",
1907 => x"a3388417",
1908 => x"08fc0670",
1909 => x"7a315556",
1910 => x"738f2483",
1911 => x"ca387380",
1912 => x"25848138",
1913 => x"8c170857",
1914 => x"76752e09",
1915 => x"8106df38",
1916 => x"8815811b",
1917 => x"70830655",
1918 => x"5b5572c9",
1919 => x"387c8306",
1920 => x"5372802e",
1921 => x"fdb838ff",
1922 => x"1df81959",
1923 => x"5d881808",
1924 => x"782eea38",
1925 => x"fdb53983",
1926 => x"1a53fc96",
1927 => x"39831470",
1928 => x"822c8171",
1929 => x"2b80d6f8",
1930 => x"08077080",
1931 => x"d6f40b84",
1932 => x"050c7610",
1933 => x"101080d6",
1934 => x"f4058811",
1935 => x"08595b5e",
1936 => x"5153fee1",
1937 => x"3980d6b8",
1938 => x"081758b0",
1939 => x"08762e81",
1940 => x"8d3880d6",
1941 => x"e808ff2e",
1942 => x"83ec3873",
1943 => x"76311880",
1944 => x"d6b80c73",
1945 => x"87067057",
1946 => x"5372802e",
1947 => x"88388873",
1948 => x"31701555",
1949 => x"5676149f",
1950 => x"ff06a080",
1951 => x"71311770",
1952 => x"547f5357",
1953 => x"5384e43f",
1954 => x"b00853b0",
1955 => x"08ff2e81",
1956 => x"a03880d6",
1957 => x"b8081670",
1958 => x"80d6b80c",
1959 => x"747580d6",
1960 => x"f40b8805",
1961 => x"0c747631",
1962 => x"18708107",
1963 => x"51555658",
1964 => x"7b80d6f4",
1965 => x"2e839c38",
1966 => x"798f2682",
1967 => x"cb38810b",
1968 => x"84150c84",
1969 => x"1508fc06",
1970 => x"707a317a",
1971 => x"72268f72",
1972 => x"25075255",
1973 => x"5372802e",
1974 => x"fcf93880",
1975 => x"db39b008",
1976 => x"9fff0653",
1977 => x"72feeb38",
1978 => x"7780d6b8",
1979 => x"0c80d6f4",
1980 => x"0b880508",
1981 => x"7b188107",
1982 => x"84120c55",
1983 => x"80d6e408",
1984 => x"78278638",
1985 => x"7780d6e4",
1986 => x"0c80d6e0",
1987 => x"087827fc",
1988 => x"ac387780",
1989 => x"d6e00c84",
1990 => x"1508fc06",
1991 => x"707a317a",
1992 => x"72268f72",
1993 => x"25075255",
1994 => x"5372802e",
1995 => x"fca53888",
1996 => x"39807454",
1997 => x"56fedb39",
1998 => x"7d5183ae",
1999 => x"3f800bb0",
2000 => x"0c8f3d0d",
2001 => x"04735380",
2002 => x"7424a938",
2003 => x"72822c81",
2004 => x"712b80d6",
2005 => x"f8080770",
2006 => x"80d6f40b",
2007 => x"84050c5d",
2008 => x"53778c18",
2009 => x"0c748818",
2010 => x"0c768819",
2011 => x"0c768c16",
2012 => x"0cf9b739",
2013 => x"83147082",
2014 => x"2c81712b",
2015 => x"80d6f808",
2016 => x"077080d6",
2017 => x"f40b8405",
2018 => x"0c5e5153",
2019 => x"d4397b7b",
2020 => x"065372fc",
2021 => x"a338841a",
2022 => x"7b105c5a",
2023 => x"f139ff1a",
2024 => x"8111515a",
2025 => x"f7b93978",
2026 => x"17798107",
2027 => x"84190c8c",
2028 => x"18088819",
2029 => x"08718c12",
2030 => x"0c88120c",
2031 => x"597080d7",
2032 => x"880c7080",
2033 => x"d7840c80",
2034 => x"d6fc0b8c",
2035 => x"120c8c11",
2036 => x"0888120c",
2037 => x"74810784",
2038 => x"120c7411",
2039 => x"75710c51",
2040 => x"53f9bd39",
2041 => x"75178411",
2042 => x"08810784",
2043 => x"120c538c",
2044 => x"17088818",
2045 => x"08718c12",
2046 => x"0c88120c",
2047 => x"587d5181",
2048 => x"e93f8817",
2049 => x"54f5cf39",
2050 => x"7284150c",
2051 => x"f41af806",
2052 => x"70841e08",
2053 => x"81060784",
2054 => x"1e0c701d",
2055 => x"545b850b",
2056 => x"84140c85",
2057 => x"0b88140c",
2058 => x"8f7b27fd",
2059 => x"cf38881c",
2060 => x"527d51ec",
2061 => x"9e3f80d6",
2062 => x"f40b8805",
2063 => x"0880d6b8",
2064 => x"085955fd",
2065 => x"b7397780",
2066 => x"d6b80c73",
2067 => x"80d6e80c",
2068 => x"fc913972",
2069 => x"84150cfd",
2070 => x"a339fc3d",
2071 => x"0d767971",
2072 => x"028c059f",
2073 => x"05335755",
2074 => x"53558372",
2075 => x"278a3874",
2076 => x"83065170",
2077 => x"802ea238",
2078 => x"ff125271",
2079 => x"ff2e9338",
2080 => x"73737081",
2081 => x"055534ff",
2082 => x"125271ff",
2083 => x"2e098106",
2084 => x"ef3874b0",
2085 => x"0c863d0d",
2086 => x"04747488",
2087 => x"2b750770",
2088 => x"71902b07",
2089 => x"5154518f",
2090 => x"7227a538",
2091 => x"72717084",
2092 => x"05530c72",
2093 => x"71708405",
2094 => x"530c7271",
2095 => x"70840553",
2096 => x"0c727170",
2097 => x"8405530c",
2098 => x"f0125271",
2099 => x"8f26dd38",
2100 => x"83722790",
2101 => x"38727170",
2102 => x"8405530c",
2103 => x"fc125271",
2104 => x"8326f238",
2105 => x"7053ff90",
2106 => x"390404fd",
2107 => x"3d0d800b",
2108 => x"80dfac0c",
2109 => x"765184ee",
2110 => x"3fb00853",
2111 => x"b008ff2e",
2112 => x"883872b0",
2113 => x"0c853d0d",
2114 => x"0480dfac",
2115 => x"08547380",
2116 => x"2ef03875",
2117 => x"74710c52",
2118 => x"72b00c85",
2119 => x"3d0d04f9",
2120 => x"3d0d797c",
2121 => x"557b548e",
2122 => x"11227090",
2123 => x"2b70902c",
2124 => x"555780cf",
2125 => x"b8085358",
2126 => x"5683f33f",
2127 => x"b0085780",
2128 => x"0bb00824",
2129 => x"933880d0",
2130 => x"1608b008",
2131 => x"0580d017",
2132 => x"0c76b00c",
2133 => x"893d0d04",
2134 => x"8c162283",
2135 => x"dfff0655",
2136 => x"748c1723",
2137 => x"76b00c89",
2138 => x"3d0d04fa",
2139 => x"3d0d788c",
2140 => x"11227088",
2141 => x"2a708106",
2142 => x"51575856",
2143 => x"74a9388c",
2144 => x"162283df",
2145 => x"ff065574",
2146 => x"8c17237a",
2147 => x"5479538e",
2148 => x"16227090",
2149 => x"2b70902c",
2150 => x"545680cf",
2151 => x"b8085256",
2152 => x"81b23f88",
2153 => x"3d0d0482",
2154 => x"5480538e",
2155 => x"16227090",
2156 => x"2b70902c",
2157 => x"545680cf",
2158 => x"b8085257",
2159 => x"82b83f8c",
2160 => x"162283df",
2161 => x"ff065574",
2162 => x"8c17237a",
2163 => x"5479538e",
2164 => x"16227090",
2165 => x"2b70902c",
2166 => x"545680cf",
2167 => x"b8085256",
2168 => x"80f23f88",
2169 => x"3d0d04f9",
2170 => x"3d0d797c",
2171 => x"557b548e",
2172 => x"11227090",
2173 => x"2b70902c",
2174 => x"555780cf",
2175 => x"b8085358",
2176 => x"5681f33f",
2177 => x"b00857b0",
2178 => x"08ff2e99",
2179 => x"388c1622",
2180 => x"a0800755",
2181 => x"748c1723",
2182 => x"b00880d0",
2183 => x"170c76b0",
2184 => x"0c893d0d",
2185 => x"048c1622",
2186 => x"83dfff06",
2187 => x"55748c17",
2188 => x"2376b00c",
2189 => x"893d0d04",
2190 => x"fe3d0d74",
2191 => x"8e112270",
2192 => x"902b7090",
2193 => x"2c555151",
2194 => x"5380cfb8",
2195 => x"0851bd3f",
2196 => x"843d0d04",
2197 => x"fb3d0d80",
2198 => x"0b80dfac",
2199 => x"0c7a5379",
2200 => x"52785182",
2201 => x"f93fb008",
2202 => x"55b008ff",
2203 => x"2e883874",
2204 => x"b00c873d",
2205 => x"0d0480df",
2206 => x"ac085675",
2207 => x"802ef038",
2208 => x"7776710c",
2209 => x"5474b00c",
2210 => x"873d0d04",
2211 => x"fd3d0d80",
2212 => x"0b80dfac",
2213 => x"0c765184",
2214 => x"c73fb008",
2215 => x"53b008ff",
2216 => x"2e883872",
2217 => x"b00c853d",
2218 => x"0d0480df",
2219 => x"ac085473",
2220 => x"802ef038",
2221 => x"7574710c",
2222 => x"5272b00c",
2223 => x"853d0d04",
2224 => x"fc3d0d80",
2225 => x"0b80dfac",
2226 => x"0c785277",
2227 => x"5186af3f",
2228 => x"b00854b0",
2229 => x"08ff2e88",
2230 => x"3873b00c",
2231 => x"863d0d04",
2232 => x"80dfac08",
2233 => x"5574802e",
2234 => x"f0387675",
2235 => x"710c5373",
2236 => x"b00c863d",
2237 => x"0d04fb3d",
2238 => x"0d800b80",
2239 => x"dfac0c7a",
2240 => x"53795278",
2241 => x"51848b3f",
2242 => x"b00855b0",
2243 => x"08ff2e88",
2244 => x"3874b00c",
2245 => x"873d0d04",
2246 => x"80dfac08",
2247 => x"5675802e",
2248 => x"f0387776",
2249 => x"710c5474",
2250 => x"b00c873d",
2251 => x"0d04fb3d",
2252 => x"0d800b80",
2253 => x"dfac0c7a",
2254 => x"53795278",
2255 => x"5182933f",
2256 => x"b00855b0",
2257 => x"08ff2e88",
2258 => x"3874b00c",
2259 => x"873d0d04",
2260 => x"80dfac08",
2261 => x"5675802e",
2262 => x"f0387776",
2263 => x"710c5474",
2264 => x"b00c873d",
2265 => x"0d04fe3d",
2266 => x"0d80dfa4",
2267 => x"0851708a",
2268 => x"3880dfb0",
2269 => x"7080dfa4",
2270 => x"0c517075",
2271 => x"125252ff",
2272 => x"537087fb",
2273 => x"80802688",
2274 => x"387080df",
2275 => x"a40c7153",
2276 => x"72b00c84",
2277 => x"3d0d04fd",
2278 => x"3d0d800b",
2279 => x"80cfa408",
2280 => x"54547281",
2281 => x"2e9b3873",
2282 => x"80dfa80c",
2283 => x"c2b83fc0",
2284 => x"cf3f80de",
2285 => x"fc528151",
2286 => x"c4e03fb0",
2287 => x"085185be",
2288 => x"3f7280df",
2289 => x"a80cc29e",
2290 => x"3fc0b53f",
2291 => x"80defc52",
2292 => x"8151c4c6",
2293 => x"3fb00851",
2294 => x"85a43f00",
2295 => x"ff39f53d",
2296 => x"0d7e6080",
2297 => x"dfa80870",
2298 => x"5b585b5b",
2299 => x"7580c238",
2300 => x"777a25a1",
2301 => x"38771b70",
2302 => x"337081ff",
2303 => x"06585859",
2304 => x"758a2e98",
2305 => x"387681ff",
2306 => x"0651c1b9",
2307 => x"3f811858",
2308 => x"797824e1",
2309 => x"3879b00c",
2310 => x"8d3d0d04",
2311 => x"8d51c1a5",
2312 => x"3f783370",
2313 => x"81ff0652",
2314 => x"57c19a3f",
2315 => x"811858e0",
2316 => x"3979557a",
2317 => x"547d5385",
2318 => x"528d3dfc",
2319 => x"0551c082",
2320 => x"3fb00856",
2321 => x"84b13f7b",
2322 => x"b0080c75",
2323 => x"b00c8d3d",
2324 => x"0d04f63d",
2325 => x"0d7d7f80",
2326 => x"dfa80870",
2327 => x"5b585a5a",
2328 => x"7580c138",
2329 => x"777925b3",
2330 => x"38c0b53f",
2331 => x"b00881ff",
2332 => x"06708d32",
2333 => x"7030709f",
2334 => x"2a515157",
2335 => x"57768a2e",
2336 => x"80c43875",
2337 => x"802ebf38",
2338 => x"771a5676",
2339 => x"76347651",
2340 => x"c0b33f81",
2341 => x"18587878",
2342 => x"24cf3877",
2343 => x"5675b00c",
2344 => x"8c3d0d04",
2345 => x"78557954",
2346 => x"7c538452",
2347 => x"8c3dfc05",
2348 => x"51ffbf8e",
2349 => x"3fb00856",
2350 => x"83bd3f7a",
2351 => x"b0080c75",
2352 => x"b00c8c3d",
2353 => x"0d04771a",
2354 => x"568a7634",
2355 => x"8118588d",
2356 => x"51ffbff1",
2357 => x"3f8a51ff",
2358 => x"bfeb3f77",
2359 => x"56ffbe39",
2360 => x"fb3d0d80",
2361 => x"dfa80870",
2362 => x"56547388",
2363 => x"3874b00c",
2364 => x"873d0d04",
2365 => x"77538352",
2366 => x"873dfc05",
2367 => x"51ffbec2",
2368 => x"3fb00854",
2369 => x"82f13f75",
2370 => x"b0080c73",
2371 => x"b00c873d",
2372 => x"0d04fa3d",
2373 => x"0d80dfa8",
2374 => x"08802ea3",
2375 => x"387a5579",
2376 => x"54785386",
2377 => x"52883dfc",
2378 => x"0551ffbe",
2379 => x"953fb008",
2380 => x"5682c43f",
2381 => x"76b0080c",
2382 => x"75b00c88",
2383 => x"3d0d0482",
2384 => x"b63f9d0b",
2385 => x"b0080cff",
2386 => x"0bb00c88",
2387 => x"3d0d04fb",
2388 => x"3d0d7779",
2389 => x"56568070",
2390 => x"54547375",
2391 => x"259f3874",
2392 => x"101010f8",
2393 => x"05527216",
2394 => x"70337074",
2395 => x"2b760781",
2396 => x"16f81656",
2397 => x"56565151",
2398 => x"747324ea",
2399 => x"3873b00c",
2400 => x"873d0d04",
2401 => x"fc3d0d76",
2402 => x"785555bc",
2403 => x"53805273",
2404 => x"51f5c73f",
2405 => x"84527451",
2406 => x"ffb53fb0",
2407 => x"08742384",
2408 => x"52841551",
2409 => x"ffa93fb0",
2410 => x"08821523",
2411 => x"84528815",
2412 => x"51ff9c3f",
2413 => x"b0088415",
2414 => x"0c84528c",
2415 => x"1551ff8f",
2416 => x"3fb00888",
2417 => x"15238452",
2418 => x"901551ff",
2419 => x"823fb008",
2420 => x"8a152384",
2421 => x"52941551",
2422 => x"fef53fb0",
2423 => x"088c1523",
2424 => x"84529815",
2425 => x"51fee83f",
2426 => x"b0088e15",
2427 => x"2388529c",
2428 => x"1551fedb",
2429 => x"3fb00890",
2430 => x"150c863d",
2431 => x"0d04e93d",
2432 => x"0d6a80df",
2433 => x"a8085757",
2434 => x"75933880",
2435 => x"c0800b84",
2436 => x"180c75ac",
2437 => x"180c75b0",
2438 => x"0c993d0d",
2439 => x"04893d70",
2440 => x"556a5455",
2441 => x"8a52993d",
2442 => x"ffbc0551",
2443 => x"ffbc933f",
2444 => x"b0087753",
2445 => x"755256fe",
2446 => x"cb3fbc3f",
2447 => x"77b0080c",
2448 => x"75b00c99",
2449 => x"3d0d04fc",
2450 => x"3d0d8154",
2451 => x"80dfa808",
2452 => x"883873b0",
2453 => x"0c863d0d",
2454 => x"04765397",
2455 => x"b952863d",
2456 => x"fc0551ff",
2457 => x"bbdc3fb0",
2458 => x"08548c3f",
2459 => x"74b0080c",
2460 => x"73b00c86",
2461 => x"3d0d0480",
2462 => x"cfb808b0",
2463 => x"0c04f73d",
2464 => x"0d7b80cf",
2465 => x"b80882c8",
2466 => x"11085a54",
2467 => x"5a77802e",
2468 => x"80da3881",
2469 => x"88188419",
2470 => x"08ff0581",
2471 => x"712b5955",
2472 => x"59807424",
2473 => x"80ea3880",
2474 => x"7424b538",
2475 => x"73822b78",
2476 => x"11880556",
2477 => x"56818019",
2478 => x"08770653",
2479 => x"72802eb6",
2480 => x"38781670",
2481 => x"08535379",
2482 => x"51740853",
2483 => x"722dff14",
2484 => x"fc17fc17",
2485 => x"79812c5a",
2486 => x"57575473",
2487 => x"8025d638",
2488 => x"77085877",
2489 => x"ffad3880",
2490 => x"cfb80853",
2491 => x"bc1308a5",
2492 => x"387951f9",
2493 => x"e63f7408",
2494 => x"53722dff",
2495 => x"14fc17fc",
2496 => x"1779812c",
2497 => x"5a575754",
2498 => x"738025ff",
2499 => x"a838d139",
2500 => x"8057ff93",
2501 => x"397251bc",
2502 => x"13085372",
2503 => x"2d7951f9",
2504 => x"ba3fff3d",
2505 => x"0d80df84",
2506 => x"0bfc0570",
2507 => x"08525270",
2508 => x"ff2e9138",
2509 => x"702dfc12",
2510 => x"70085252",
2511 => x"70ff2e09",
2512 => x"8106f138",
2513 => x"833d0d04",
2514 => x"04ffbc85",
2515 => x"3f040000",
2516 => x"00ffffff",
2517 => x"ff00ffff",
2518 => x"ffff00ff",
2519 => x"ffffff00",
2520 => x"00000040",
2521 => x"30313233",
2522 => x"34353637",
2523 => x"38396162",
2524 => x"63646566",
2525 => x"00000000",
2526 => x"2d2d0000",
2527 => x"6c6f6f70",
2528 => x"00000000",
2529 => x"636e743a",
2530 => x"20000000",
2531 => x"0a000000",
2532 => x"43000000",
2533 => x"64756d6d",
2534 => x"792e6578",
2535 => x"65000000",
2536 => x"00000000",
2537 => x"00000000",
2538 => x"00000000",
2539 => x"00002f8c",
2540 => x"00000000",
2541 => x"00002764",
2542 => x"000027bc",
2543 => x"00000000",
2544 => x"00002a24",
2545 => x"00002a80",
2546 => x"00002adc",
2547 => x"00000000",
2548 => x"00000000",
2549 => x"00000000",
2550 => x"00000000",
2551 => x"00000000",
2552 => x"00000000",
2553 => x"00000000",
2554 => x"00000000",
2555 => x"00000000",
2556 => x"00002790",
2557 => x"00000000",
2558 => x"00000000",
2559 => x"00000000",
2560 => x"00000000",
2561 => x"00000000",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"00000000",
2568 => x"00000000",
2569 => x"00000000",
2570 => x"00000000",
2571 => x"00000000",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000001",
2586 => x"330eabcd",
2587 => x"1234e66d",
2588 => x"deec0005",
2589 => x"000b0000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000000",
2597 => x"00000000",
2598 => x"00000000",
2599 => x"00000000",
2600 => x"00000000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"ffffffff",
2779 => x"00000000",
2780 => x"00020000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00002b74",
2784 => x"00002b74",
2785 => x"00002b7c",
2786 => x"00002b7c",
2787 => x"00002b84",
2788 => x"00002b84",
2789 => x"00002b8c",
2790 => x"00002b8c",
2791 => x"00002b94",
2792 => x"00002b94",
2793 => x"00002b9c",
2794 => x"00002b9c",
2795 => x"00002ba4",
2796 => x"00002ba4",
2797 => x"00002bac",
2798 => x"00002bac",
2799 => x"00002bb4",
2800 => x"00002bb4",
2801 => x"00002bbc",
2802 => x"00002bbc",
2803 => x"00002bc4",
2804 => x"00002bc4",
2805 => x"00002bcc",
2806 => x"00002bcc",
2807 => x"00002bd4",
2808 => x"00002bd4",
2809 => x"00002bdc",
2810 => x"00002bdc",
2811 => x"00002be4",
2812 => x"00002be4",
2813 => x"00002bec",
2814 => x"00002bec",
2815 => x"00002bf4",
2816 => x"00002bf4",
2817 => x"00002bfc",
2818 => x"00002bfc",
2819 => x"00002c04",
2820 => x"00002c04",
2821 => x"00002c0c",
2822 => x"00002c0c",
2823 => x"00002c14",
2824 => x"00002c14",
2825 => x"00002c1c",
2826 => x"00002c1c",
2827 => x"00002c24",
2828 => x"00002c24",
2829 => x"00002c2c",
2830 => x"00002c2c",
2831 => x"00002c34",
2832 => x"00002c34",
2833 => x"00002c3c",
2834 => x"00002c3c",
2835 => x"00002c44",
2836 => x"00002c44",
2837 => x"00002c4c",
2838 => x"00002c4c",
2839 => x"00002c54",
2840 => x"00002c54",
2841 => x"00002c5c",
2842 => x"00002c5c",
2843 => x"00002c64",
2844 => x"00002c64",
2845 => x"00002c6c",
2846 => x"00002c6c",
2847 => x"00002c74",
2848 => x"00002c74",
2849 => x"00002c7c",
2850 => x"00002c7c",
2851 => x"00002c84",
2852 => x"00002c84",
2853 => x"00002c8c",
2854 => x"00002c8c",
2855 => x"00002c94",
2856 => x"00002c94",
2857 => x"00002c9c",
2858 => x"00002c9c",
2859 => x"00002ca4",
2860 => x"00002ca4",
2861 => x"00002cac",
2862 => x"00002cac",
2863 => x"00002cb4",
2864 => x"00002cb4",
2865 => x"00002cbc",
2866 => x"00002cbc",
2867 => x"00002cc4",
2868 => x"00002cc4",
2869 => x"00002ccc",
2870 => x"00002ccc",
2871 => x"00002cd4",
2872 => x"00002cd4",
2873 => x"00002cdc",
2874 => x"00002cdc",
2875 => x"00002ce4",
2876 => x"00002ce4",
2877 => x"00002cec",
2878 => x"00002cec",
2879 => x"00002cf4",
2880 => x"00002cf4",
2881 => x"00002cfc",
2882 => x"00002cfc",
2883 => x"00002d04",
2884 => x"00002d04",
2885 => x"00002d0c",
2886 => x"00002d0c",
2887 => x"00002d14",
2888 => x"00002d14",
2889 => x"00002d1c",
2890 => x"00002d1c",
2891 => x"00002d24",
2892 => x"00002d24",
2893 => x"00002d2c",
2894 => x"00002d2c",
2895 => x"00002d34",
2896 => x"00002d34",
2897 => x"00002d3c",
2898 => x"00002d3c",
2899 => x"00002d44",
2900 => x"00002d44",
2901 => x"00002d4c",
2902 => x"00002d4c",
2903 => x"00002d54",
2904 => x"00002d54",
2905 => x"00002d5c",
2906 => x"00002d5c",
2907 => x"00002d64",
2908 => x"00002d64",
2909 => x"00002d6c",
2910 => x"00002d6c",
2911 => x"00002d74",
2912 => x"00002d74",
2913 => x"00002d7c",
2914 => x"00002d7c",
2915 => x"00002d84",
2916 => x"00002d84",
2917 => x"00002d8c",
2918 => x"00002d8c",
2919 => x"00002d94",
2920 => x"00002d94",
2921 => x"00002d9c",
2922 => x"00002d9c",
2923 => x"00002da4",
2924 => x"00002da4",
2925 => x"00002dac",
2926 => x"00002dac",
2927 => x"00002db4",
2928 => x"00002db4",
2929 => x"00002dbc",
2930 => x"00002dbc",
2931 => x"00002dc4",
2932 => x"00002dc4",
2933 => x"00002dcc",
2934 => x"00002dcc",
2935 => x"00002dd4",
2936 => x"00002dd4",
2937 => x"00002ddc",
2938 => x"00002ddc",
2939 => x"00002de4",
2940 => x"00002de4",
2941 => x"00002dec",
2942 => x"00002dec",
2943 => x"00002df4",
2944 => x"00002df4",
2945 => x"00002dfc",
2946 => x"00002dfc",
2947 => x"00002e04",
2948 => x"00002e04",
2949 => x"00002e0c",
2950 => x"00002e0c",
2951 => x"00002e14",
2952 => x"00002e14",
2953 => x"00002e1c",
2954 => x"00002e1c",
2955 => x"00002e24",
2956 => x"00002e24",
2957 => x"00002e2c",
2958 => x"00002e2c",
2959 => x"00002e34",
2960 => x"00002e34",
2961 => x"00002e3c",
2962 => x"00002e3c",
2963 => x"00002e44",
2964 => x"00002e44",
2965 => x"00002e4c",
2966 => x"00002e4c",
2967 => x"00002e54",
2968 => x"00002e54",
2969 => x"00002e5c",
2970 => x"00002e5c",
2971 => x"00002e64",
2972 => x"00002e64",
2973 => x"00002e6c",
2974 => x"00002e6c",
2975 => x"00002e74",
2976 => x"00002e74",
2977 => x"00002e7c",
2978 => x"00002e7c",
2979 => x"00002e84",
2980 => x"00002e84",
2981 => x"00002e8c",
2982 => x"00002e8c",
2983 => x"00002e94",
2984 => x"00002e94",
2985 => x"00002e9c",
2986 => x"00002e9c",
2987 => x"00002ea4",
2988 => x"00002ea4",
2989 => x"00002eac",
2990 => x"00002eac",
2991 => x"00002eb4",
2992 => x"00002eb4",
2993 => x"00002ebc",
2994 => x"00002ebc",
2995 => x"00002ec4",
2996 => x"00002ec4",
2997 => x"00002ecc",
2998 => x"00002ecc",
2999 => x"00002ed4",
3000 => x"00002ed4",
3001 => x"00002edc",
3002 => x"00002edc",
3003 => x"00002ee4",
3004 => x"00002ee4",
3005 => x"00002eec",
3006 => x"00002eec",
3007 => x"00002ef4",
3008 => x"00002ef4",
3009 => x"00002efc",
3010 => x"00002efc",
3011 => x"00002f04",
3012 => x"00002f04",
3013 => x"00002f0c",
3014 => x"00002f0c",
3015 => x"00002f14",
3016 => x"00002f14",
3017 => x"00002f1c",
3018 => x"00002f1c",
3019 => x"00002f24",
3020 => x"00002f24",
3021 => x"00002f2c",
3022 => x"00002f2c",
3023 => x"00002f34",
3024 => x"00002f34",
3025 => x"00002f3c",
3026 => x"00002f3c",
3027 => x"00002f44",
3028 => x"00002f44",
3029 => x"00002f4c",
3030 => x"00002f4c",
3031 => x"00002f54",
3032 => x"00002f54",
3033 => x"00002f5c",
3034 => x"00002f5c",
3035 => x"00002f64",
3036 => x"00002f64",
3037 => x"00002f6c",
3038 => x"00002f6c",
3039 => x"00002794",
3040 => x"ffffffff",
3041 => x"00000000",
3042 => x"ffffffff",
3043 => x"00000000",
others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

